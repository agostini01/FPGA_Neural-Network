-------------------------------------------------------
-- Design Name : User Pakage
-- File Name   : neural_net_pkg.vhd
-- Function    : 
-- Coder       : Agostini, N. & Barbosa, F.
-------------------------------------------------------
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;

	use work.fixed_float_types.all; -- ieee_proposed for VHDL-93 version
	use work.fixed_pkg.all; -- ieee_proposed for compatibility version

package NN_PKG is


			constant INPUT_PERCEPTRONS 	: natural := 13;
			constant HIDDEN_PERCEPTRONS 	: natural := 4;
			constant OUT_PERCEPTRONS 		: natural := 3;
			
			constant F_U_SIZE : integer :=11;
			constant F_L_SIZE : integer :=-4;
		--	constant FIX_SIZE 	: sfixed := to_sfixed(6.5 ,5,-2);
			type INT_ARRAY is array (natural range <>) of natural;
			
			subtype S_SFIXED is sfixed(F_U_SIZE downto F_L_SIZE);
			type FIX_ARRAY is array (natural range <>) of S_SFIXED;
			
			subtype IN_FIX_ARRAY is FIX_ARRAY  (0 to (INPUT_PERCEPTRONS-1));
			subtype HID_FIX_ARRAY is FIX_ARRAY  (0 to (HIDDEN_PERCEPTRONS-1));
			subtype OUT_FIX_ARRAY is FIX_ARRAY  (0 to (OUT_PERCEPTRONS-1));
			type FIX_ARRAY_2D is array (natural range <>) of FIX_ARRAY(open);
			type FIX_ARRAY_3D is array (natural range <>) of FIX_ARRAY_2D;


			
			
			type T_WINE_DATASET is array (0 to 177, 0 to 13) of S_SFIXED;

			


end;

package body NN_PKG is
	
	-- biases and weights for input layer
	constant wine_dataset_init_input_layer : FIX_ARRAY_2D(0 to 12) := (
	
	-- biases and weights for hidden layer
		(to_sfixed(1,11,-4),to_sfixed(0,11,-4)),
		(to_sfixed(1,11,-4),to_sfixed(0,11,-4)),
		(to_sfixed(1,11,-4),to_sfixed(0,11,-4)),
		(to_sfixed(1,11,-4),to_sfixed(0,11,-4)),
		(to_sfixed(1,11,-4),to_sfixed(0,11,-4)),
		(to_sfixed(1,11,-4),to_sfixed(0,11,-4)),
		(to_sfixed(1,11,-4),to_sfixed(0,11,-4)),
		(to_sfixed(1,11,-4),to_sfixed(0,11,-4)),
		(to_sfixed(1,11,-4),to_sfixed(0,11,-4)),
		(to_sfixed(1,11,-4),to_sfixed(0,11,-4)),
		(to_sfixed(1,11,-4),to_sfixed(0,11,-4)),
		(to_sfixed(1,11,-4),to_sfixed(0,11,-4)),
		(to_sfixed(1,11,-4),to_sfixed(0,11,-4))
	);

	constant wine_dataset_init_hidden_layer : FIX_ARRAY_2D(0 to 2) := (
	
	-- biases and weights for output layer
		(to_sfixed(-0.2944,11,-4),to_sfixed(-0.1762,11,-4),to_sfixed(0.0424,11,-4),to_sfixed(0.4687,11,-4),to_sfixed(-0.5961,11,-4),to_sfixed(-0.7336,11,-4),to_sfixed(0.0010,11,-4),to_sfixed(-0.4148,11,-4),to_sfixed(-0.2067,11,-4),to_sfixed(0.1213,11,-4),to_sfixed(0.1815,11,-4),to_sfixed(-0.3707,11,-4),to_sfixed(0.1376,11,-4),to_sfixed(2.1061,11,-4)),
		(to_sfixed(-1.9218,11,-4),to_sfixed(-0.8591,11,-4),to_sfixed(-2.2805,11,-4),to_sfixed(2.3456,11,-4),to_sfixed(-0.1239,11,-4),to_sfixed(-0.0335,11,-4),to_sfixed(-0.6953,11,-4),to_sfixed(0.0853,11,-4),to_sfixed(-0.0385,11,-4),to_sfixed(-0.4995,11,-4),to_sfixed(0.6088,11,-4),to_sfixed(-1.4969,11,-4),to_sfixed(-2.6136,11,-4),to_sfixed(-0.4546,11,-4)),
		(to_sfixed(-0.3840,11,-4),to_sfixed(-0.6723,11,-4),to_sfixed(-0.5043,11,-4),to_sfixed(-0.3566,11,-4),to_sfixed(-0.0082,11,-4),to_sfixed(-0.6894,11,-4),to_sfixed(2.8733,11,-4),to_sfixed(0.7266,11,-4),to_sfixed(1.0385,11,-4),to_sfixed(-2.8766,11,-4),to_sfixed(1.5652,11,-4),to_sfixed(1.8564,11,-4),to_sfixed(-0.3278,11,-4),to_sfixed(1.9498,11,-4))
	);

	constant wine_dataset_init_output_layer : FIX_ARRAY_2D(0 to 2) := (
	
	-- biases and weights matrix
		(to_sfixed(-1.9038,11,-4),to_sfixed(-4.1782,11,-4),to_sfixed(1.3133,11,-4),to_sfixed(0.4581,11,-4)),
		(to_sfixed(-1.7035,11,-4),to_sfixed(4.1581,11,-4),to_sfixed(3.9893,11,-4),to_sfixed(-2.2319,11,-4)),
		(to_sfixed(0.2439,11,-4),to_sfixed(0.0295,11,-4),to_sfixed(-4.1666,11,-4),to_sfixed(-0.3156,11,-4))
	);
	
	constant wine_dataset_init_layer_matrix : FIX_ARRAY_3D(0 to 2) := (
	
	-- wine dataset (https://archive.ics.uci.edu/ml/datasets/Wine)
		(wine_dataset_init_input_layer), 
		(wine_dataset_init_hidden_layer), 
		(wine_dataset_init_output_layer)
	);

	constant wine_dataset : T_WINE_DATASET := (

		(
		to_sfixed(1,11,-4),
		to_sfixed(14.23,11,-4),
		to_sfixed(1.71,11,-4),
		to_sfixed(2.43,11,-4),
		to_sfixed(15.6,11,-4),
		to_sfixed(127.0,11,-4),
		to_sfixed(2.8,11,-4),
		to_sfixed(3.06,11,-4),
		to_sfixed(0.28,11,-4),
		to_sfixed(2.29,11,-4),
		to_sfixed(5.64,11,-4),
		to_sfixed(1.04,11,-4),
		to_sfixed(3.92,11,-4),
		to_sfixed(1065.0,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.2,11,-4),
		to_sfixed(1.78,11,-4),
		to_sfixed(2.14,11,-4),
		to_sfixed(11.2,11,-4),
		to_sfixed(100,11,-4),
		to_sfixed(2.65,11,-4),
		to_sfixed(2.76,11,-4),
		to_sfixed(0.26,11,-4),
		to_sfixed(1.28,11,-4),
		to_sfixed(4.38,11,-4),
		to_sfixed(1.05,11,-4),
		to_sfixed(3.4,11,-4),
		to_sfixed(1050,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.16,11,-4),
		to_sfixed(2.36,11,-4),
		to_sfixed(2.67,11,-4),
		to_sfixed(18.6,11,-4),
		to_sfixed(101,11,-4),
		to_sfixed(2.8,11,-4),
		to_sfixed(3.24,11,-4),
		to_sfixed(0.3,11,-4),
		to_sfixed(2.81,11,-4),
		to_sfixed(5.68,11,-4),
		to_sfixed(1.03,11,-4),
		to_sfixed(3.17,11,-4),
		to_sfixed(1185,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(14.37,11,-4),
		to_sfixed(1.95,11,-4),
		to_sfixed(2.50,11,-4),
		to_sfixed(16.8,11,-4),
		to_sfixed(113,11,-4),
		to_sfixed(3.85,11,-4),
		to_sfixed(3.49,11,-4),
		to_sfixed(0.24,11,-4),
		to_sfixed(2.18,11,-4),
		to_sfixed(7.8,11,-4),
		to_sfixed(0.86,11,-4),
		to_sfixed(3.45,11,-4),
		to_sfixed(1480,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.24,11,-4),
		to_sfixed(2.59,11,-4),
		to_sfixed(2.87,11,-4),
		to_sfixed(21,11,-4),
		to_sfixed(118,11,-4),
		to_sfixed(2.8,11,-4),
		to_sfixed(2.69,11,-4),
		to_sfixed(0.39,11,-4),
		to_sfixed(1.82,11,-4),
		to_sfixed(4.32,11,-4),
		to_sfixed(1.04,11,-4),
		to_sfixed(2.93,11,-4),
		to_sfixed(735,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(14.2,11,-4),
		to_sfixed(1.76,11,-4),
		to_sfixed(2.45,11,-4),
		to_sfixed(15.2,11,-4),
		to_sfixed(112,11,-4),
		to_sfixed(3.27,11,-4),
		to_sfixed(3.39,11,-4),
		to_sfixed(0.34,11,-4),
		to_sfixed(1.97,11,-4),
		to_sfixed(6.75,11,-4),
		to_sfixed(1.05,11,-4),
		to_sfixed(2.85,11,-4),
		to_sfixed(1450,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(14.39,11,-4),
		to_sfixed(1.87,11,-4),
		to_sfixed(2.45,11,-4),
		to_sfixed(14.6,11,-4),
		to_sfixed(96,11,-4),
		to_sfixed(2.5,11,-4),
		to_sfixed(2.52,11,-4),
		to_sfixed(0.3,11,-4),
		to_sfixed(1.98,11,-4),
		to_sfixed(5.25,11,-4),
		to_sfixed(1.02,11,-4),
		to_sfixed(3.58,11,-4),
		to_sfixed(1290,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(14.06,11,-4),
		to_sfixed(2.15,11,-4),
		to_sfixed(2.61,11,-4),
		to_sfixed(17.6,11,-4),
		to_sfixed(121,11,-4),
		to_sfixed(2.6,11,-4),
		to_sfixed(2.51,11,-4),
		to_sfixed(0.31,11,-4),
		to_sfixed(1.25,11,-4),
		to_sfixed(5.05,11,-4),
		to_sfixed(1.06,11,-4),
		to_sfixed(3.58,11,-4),
		to_sfixed(1295,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(14.83,11,-4),
		to_sfixed(1.64,11,-4),
		to_sfixed(2.17,11,-4),
		to_sfixed(14,11,-4),
		to_sfixed(97,11,-4),
		to_sfixed(2.8,11,-4),
		to_sfixed(2.98,11,-4),
		to_sfixed(0.29,11,-4),
		to_sfixed(1.98,11,-4),
		to_sfixed(5.2,11,-4),
		to_sfixed(1.08,11,-4),
		to_sfixed(2.85,11,-4),
		to_sfixed(1045,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.86,11,-4),
		to_sfixed(1.35,11,-4),
		to_sfixed(2.27,11,-4),
		to_sfixed(16,11,-4),
		to_sfixed(98,11,-4),
		to_sfixed(2.98,11,-4),
		to_sfixed(3.15,11,-4),
		to_sfixed(0.22,11,-4),
		to_sfixed(1.85,11,-4),
		to_sfixed(7.22,11,-4),
		to_sfixed(1.01,11,-4),
		to_sfixed(3.55,11,-4),
		to_sfixed(1045,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(14.1,11,-4),
		to_sfixed(2.16,11,-4),
		to_sfixed(2.30,11,-4),
		to_sfixed(18,11,-4),
		to_sfixed(105,11,-4),
		to_sfixed(2.95,11,-4),
		to_sfixed(3.32,11,-4),
		to_sfixed(0.22,11,-4),
		to_sfixed(2.38,11,-4),
		to_sfixed(5.75,11,-4),
		to_sfixed(1.25,11,-4),
		to_sfixed(3.17,11,-4),
		to_sfixed(1510,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(14.12,11,-4),
		to_sfixed(1.48,11,-4),
		to_sfixed(2.32,11,-4),
		to_sfixed(16.8,11,-4),
		to_sfixed(95,11,-4),
		to_sfixed(2.2,11,-4),
		to_sfixed(2.43,11,-4),
		to_sfixed(0.26,11,-4),
		to_sfixed(1.57,11,-4),
		to_sfixed(5,11,-4),
		to_sfixed(1.17,11,-4),
		to_sfixed(2.82,11,-4),
		to_sfixed(1280,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.75,11,-4),
		to_sfixed(1.73,11,-4),
		to_sfixed(2.41,11,-4),
		to_sfixed(16,11,-4),
		to_sfixed(89,11,-4),
		to_sfixed(2.6,11,-4),
		to_sfixed(2.76,11,-4),
		to_sfixed(0.29,11,-4),
		to_sfixed(1.81,11,-4),
		to_sfixed(5.6,11,-4),
		to_sfixed(1.15,11,-4),
		to_sfixed(2.9,11,-4),
		to_sfixed(1320,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(14.75,11,-4),
		to_sfixed(1.73,11,-4),
		to_sfixed(2.39,11,-4),
		to_sfixed(11.4,11,-4),
		to_sfixed(91,11,-4),
		to_sfixed(3.1,11,-4),
		to_sfixed(3.69,11,-4),
		to_sfixed(0.43,11,-4),
		to_sfixed(2.81,11,-4),
		to_sfixed(5.4,11,-4),
		to_sfixed(1.25,11,-4),
		to_sfixed(2.73,11,-4),
		to_sfixed(1150,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(14.38,11,-4),
		to_sfixed(1.87,11,-4),
		to_sfixed(2.38,11,-4),
		to_sfixed(12,11,-4),
		to_sfixed(102,11,-4),
		to_sfixed(3.3,11,-4),
		to_sfixed(3.64,11,-4),
		to_sfixed(0.29,11,-4),
		to_sfixed(2.96,11,-4),
		to_sfixed(7.5,11,-4),
		to_sfixed(1.2,11,-4),
		to_sfixed(3,11,-4),
		to_sfixed(1547,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.63,11,-4),
		to_sfixed(1.81,11,-4),
		to_sfixed(2.70,11,-4),
		to_sfixed(17.2,11,-4),
		to_sfixed(112,11,-4),
		to_sfixed(2.85,11,-4),
		to_sfixed(2.91,11,-4),
		to_sfixed(0.3,11,-4),
		to_sfixed(1.46,11,-4),
		to_sfixed(7.3,11,-4),
		to_sfixed(1.28,11,-4),
		to_sfixed(2.88,11,-4),
		to_sfixed(1310,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(14.3,11,-4),
		to_sfixed(1.92,11,-4),
		to_sfixed(2.72,11,-4),
		to_sfixed(20,11,-4),
		to_sfixed(120,11,-4),
		to_sfixed(2.8,11,-4),
		to_sfixed(3.14,11,-4),
		to_sfixed(0.33,11,-4),
		to_sfixed(1.97,11,-4),
		to_sfixed(6.2,11,-4),
		to_sfixed(1.07,11,-4),
		to_sfixed(2.65,11,-4),
		to_sfixed(1280,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.83,11,-4),
		to_sfixed(1.57,11,-4),
		to_sfixed(2.62,11,-4),
		to_sfixed(20,11,-4),
		to_sfixed(115,11,-4),
		to_sfixed(2.95,11,-4),
		to_sfixed(3.4,11,-4),
		to_sfixed(0.4,11,-4),
		to_sfixed(1.72,11,-4),
		to_sfixed(6.6,11,-4),
		to_sfixed(1.13,11,-4),
		to_sfixed(2.57,11,-4),
		to_sfixed(1130,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(14.19,11,-4),
		to_sfixed(1.59,11,-4),
		to_sfixed(2.48,11,-4),
		to_sfixed(16.5,11,-4),
		to_sfixed(108,11,-4),
		to_sfixed(3.3,11,-4),
		to_sfixed(3.93,11,-4),
		to_sfixed(0.32,11,-4),
		to_sfixed(1.86,11,-4),
		to_sfixed(8.7,11,-4),
		to_sfixed(1.23,11,-4),
		to_sfixed(2.82,11,-4),
		to_sfixed(1680,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.64,11,-4),
		to_sfixed(3.10,11,-4),
		to_sfixed(2.56,11,-4),
		to_sfixed(15.2,11,-4),
		to_sfixed(116,11,-4),
		to_sfixed(2.7,11,-4),
		to_sfixed(3.03,11,-4),
		to_sfixed(0.17,11,-4),
		to_sfixed(1.66,11,-4),
		to_sfixed(5.1,11,-4),
		to_sfixed(0.96,11,-4),
		to_sfixed(3.36,11,-4),
		to_sfixed(845,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(14.06,11,-4),
		to_sfixed(1.63,11,-4),
		to_sfixed(2.28,11,-4),
		to_sfixed(16,11,-4),
		to_sfixed(126,11,-4),
		to_sfixed(3,11,-4),
		to_sfixed(3.17,11,-4),
		to_sfixed(0.24,11,-4),
		to_sfixed(2.1,11,-4),
		to_sfixed(5.65,11,-4),
		to_sfixed(1.09,11,-4),
		to_sfixed(3.71,11,-4),
		to_sfixed(780,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(12.93,11,-4),
		to_sfixed(3.80,11,-4),
		to_sfixed(2.65,11,-4),
		to_sfixed(18.6,11,-4),
		to_sfixed(102,11,-4),
		to_sfixed(2.41,11,-4),
		to_sfixed(2.41,11,-4),
		to_sfixed(0.25,11,-4),
		to_sfixed(1.98,11,-4),
		to_sfixed(4.5,11,-4),
		to_sfixed(1.03,11,-4),
		to_sfixed(3.52,11,-4),
		to_sfixed(770,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.71,11,-4),
		to_sfixed(1.86,11,-4),
		to_sfixed(2.36,11,-4),
		to_sfixed(16.6,11,-4),
		to_sfixed(101,11,-4),
		to_sfixed(2.61,11,-4),
		to_sfixed(2.88,11,-4),
		to_sfixed(0.27,11,-4),
		to_sfixed(1.69,11,-4),
		to_sfixed(3.8,11,-4),
		to_sfixed(1.11,11,-4),
		to_sfixed(4,11,-4),
		to_sfixed(1035,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(12.85,11,-4),
		to_sfixed(1.60,11,-4),
		to_sfixed(2.52,11,-4),
		to_sfixed(17.8,11,-4),
		to_sfixed(95,11,-4),
		to_sfixed(2.48,11,-4),
		to_sfixed(2.37,11,-4),
		to_sfixed(0.26,11,-4),
		to_sfixed(1.46,11,-4),
		to_sfixed(3.93,11,-4),
		to_sfixed(1.09,11,-4),
		to_sfixed(3.63,11,-4),
		to_sfixed(1015,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.5,11,-4),
		to_sfixed(1.81,11,-4),
		to_sfixed(2.61,11,-4),
		to_sfixed(20,11,-4),
		to_sfixed(96,11,-4),
		to_sfixed(2.53,11,-4),
		to_sfixed(2.61,11,-4),
		to_sfixed(0.28,11,-4),
		to_sfixed(1.66,11,-4),
		to_sfixed(3.52,11,-4),
		to_sfixed(1.12,11,-4),
		to_sfixed(3.82,11,-4),
		to_sfixed(845,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.05,11,-4),
		to_sfixed(2.05,11,-4),
		to_sfixed(3.22,11,-4),
		to_sfixed(25,11,-4),
		to_sfixed(124,11,-4),
		to_sfixed(2.63,11,-4),
		to_sfixed(2.68,11,-4),
		to_sfixed(0.47,11,-4),
		to_sfixed(1.92,11,-4),
		to_sfixed(3.58,11,-4),
		to_sfixed(1.13,11,-4),
		to_sfixed(3.2,11,-4),
		to_sfixed(830,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.39,11,-4),
		to_sfixed(1.77,11,-4),
		to_sfixed(2.62,11,-4),
		to_sfixed(16.1,11,-4),
		to_sfixed(93,11,-4),
		to_sfixed(2.85,11,-4),
		to_sfixed(2.94,11,-4),
		to_sfixed(0.34,11,-4),
		to_sfixed(1.45,11,-4),
		to_sfixed(4.8,11,-4),
		to_sfixed(0.92,11,-4),
		to_sfixed(3.22,11,-4),
		to_sfixed(1195,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.3,11,-4),
		to_sfixed(1.72,11,-4),
		to_sfixed(2.14,11,-4),
		to_sfixed(17,11,-4),
		to_sfixed(94,11,-4),
		to_sfixed(2.4,11,-4),
		to_sfixed(2.19,11,-4),
		to_sfixed(0.27,11,-4),
		to_sfixed(1.35,11,-4),
		to_sfixed(3.95,11,-4),
		to_sfixed(1.02,11,-4),
		to_sfixed(2.77,11,-4),
		to_sfixed(1285,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.87,11,-4),
		to_sfixed(1.90,11,-4),
		to_sfixed(2.80,11,-4),
		to_sfixed(19.4,11,-4),
		to_sfixed(107,11,-4),
		to_sfixed(2.95,11,-4),
		to_sfixed(2.97,11,-4),
		to_sfixed(0.37,11,-4),
		to_sfixed(1.76,11,-4),
		to_sfixed(4.5,11,-4),
		to_sfixed(1.25,11,-4),
		to_sfixed(3.4,11,-4),
		to_sfixed(915,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(14.02,11,-4),
		to_sfixed(1.68,11,-4),
		to_sfixed(2.21,11,-4),
		to_sfixed(16,11,-4),
		to_sfixed(96,11,-4),
		to_sfixed(2.65,11,-4),
		to_sfixed(2.33,11,-4),
		to_sfixed(0.26,11,-4),
		to_sfixed(1.98,11,-4),
		to_sfixed(4.7,11,-4),
		to_sfixed(1.04,11,-4),
		to_sfixed(3.59,11,-4),
		to_sfixed(1035,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.73,11,-4),
		to_sfixed(1.50,11,-4),
		to_sfixed(2.70,11,-4),
		to_sfixed(22.5,11,-4),
		to_sfixed(101,11,-4),
		to_sfixed(3,11,-4),
		to_sfixed(3.25,11,-4),
		to_sfixed(0.29,11,-4),
		to_sfixed(2.38,11,-4),
		to_sfixed(5.7,11,-4),
		to_sfixed(1.19,11,-4),
		to_sfixed(2.71,11,-4),
		to_sfixed(1285,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.58,11,-4),
		to_sfixed(1.66,11,-4),
		to_sfixed(2.36,11,-4),
		to_sfixed(19.1,11,-4),
		to_sfixed(106,11,-4),
		to_sfixed(2.86,11,-4),
		to_sfixed(3.19,11,-4),
		to_sfixed(0.22,11,-4),
		to_sfixed(1.95,11,-4),
		to_sfixed(6.9,11,-4),
		to_sfixed(1.09,11,-4),
		to_sfixed(2.88,11,-4),
		to_sfixed(1515,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.68,11,-4),
		to_sfixed(1.83,11,-4),
		to_sfixed(2.36,11,-4),
		to_sfixed(17.2,11,-4),
		to_sfixed(104,11,-4),
		to_sfixed(2.42,11,-4),
		to_sfixed(2.69,11,-4),
		to_sfixed(0.42,11,-4),
		to_sfixed(1.97,11,-4),
		to_sfixed(3.84,11,-4),
		to_sfixed(1.23,11,-4),
		to_sfixed(2.87,11,-4),
		to_sfixed(990,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.76,11,-4),
		to_sfixed(1.53,11,-4),
		to_sfixed(2.70,11,-4),
		to_sfixed(19.5,11,-4),
		to_sfixed(132,11,-4),
		to_sfixed(2.95,11,-4),
		to_sfixed(2.74,11,-4),
		to_sfixed(0.5,11,-4),
		to_sfixed(1.35,11,-4),
		to_sfixed(5.4,11,-4),
		to_sfixed(1.25,11,-4),
		to_sfixed(3,11,-4),
		to_sfixed(1235,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.51,11,-4),
		to_sfixed(1.80,11,-4),
		to_sfixed(2.65,11,-4),
		to_sfixed(19,11,-4),
		to_sfixed(110,11,-4),
		to_sfixed(2.35,11,-4),
		to_sfixed(2.53,11,-4),
		to_sfixed(0.29,11,-4),
		to_sfixed(1.54,11,-4),
		to_sfixed(4.2,11,-4),
		to_sfixed(1.1,11,-4),
		to_sfixed(2.87,11,-4),
		to_sfixed(1095,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.48,11,-4),
		to_sfixed(1.81,11,-4),
		to_sfixed(2.41,11,-4),
		to_sfixed(20.5,11,-4),
		to_sfixed(100,11,-4),
		to_sfixed(2.7,11,-4),
		to_sfixed(2.98,11,-4),
		to_sfixed(0.26,11,-4),
		to_sfixed(1.86,11,-4),
		to_sfixed(5.1,11,-4),
		to_sfixed(1.04,11,-4),
		to_sfixed(3.47,11,-4),
		to_sfixed(920,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.28,11,-4),
		to_sfixed(1.64,11,-4),
		to_sfixed(2.84,11,-4),
		to_sfixed(15.5,11,-4),
		to_sfixed(110,11,-4),
		to_sfixed(2.6,11,-4),
		to_sfixed(2.68,11,-4),
		to_sfixed(0.34,11,-4),
		to_sfixed(1.36,11,-4),
		to_sfixed(4.6,11,-4),
		to_sfixed(1.09,11,-4),
		to_sfixed(2.78,11,-4),
		to_sfixed(880,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.05,11,-4),
		to_sfixed(1.65,11,-4),
		to_sfixed(2.55,11,-4),
		to_sfixed(18,11,-4),
		to_sfixed(98,11,-4),
		to_sfixed(2.45,11,-4),
		to_sfixed(2.43,11,-4),
		to_sfixed(0.29,11,-4),
		to_sfixed(1.44,11,-4),
		to_sfixed(4.25,11,-4),
		to_sfixed(1.12,11,-4),
		to_sfixed(2.51,11,-4),
		to_sfixed(1105,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.07,11,-4),
		to_sfixed(1.50,11,-4),
		to_sfixed(2.10,11,-4),
		to_sfixed(15.5,11,-4),
		to_sfixed(98,11,-4),
		to_sfixed(2.4,11,-4),
		to_sfixed(2.64,11,-4),
		to_sfixed(0.28,11,-4),
		to_sfixed(1.37,11,-4),
		to_sfixed(3.7,11,-4),
		to_sfixed(1.18,11,-4),
		to_sfixed(2.69,11,-4),
		to_sfixed(1020,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(14.22,11,-4),
		to_sfixed(3.99,11,-4),
		to_sfixed(2.51,11,-4),
		to_sfixed(13.2,11,-4),
		to_sfixed(128,11,-4),
		to_sfixed(3,11,-4),
		to_sfixed(3.04,11,-4),
		to_sfixed(0.2,11,-4),
		to_sfixed(2.08,11,-4),
		to_sfixed(5.1,11,-4),
		to_sfixed(0.89,11,-4),
		to_sfixed(3.53,11,-4),
		to_sfixed(760,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.56,11,-4),
		to_sfixed(1.71,11,-4),
		to_sfixed(2.31,11,-4),
		to_sfixed(16.2,11,-4),
		to_sfixed(117,11,-4),
		to_sfixed(3.15,11,-4),
		to_sfixed(3.29,11,-4),
		to_sfixed(0.34,11,-4),
		to_sfixed(2.34,11,-4),
		to_sfixed(6.13,11,-4),
		to_sfixed(0.95,11,-4),
		to_sfixed(3.38,11,-4),
		to_sfixed(795,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.41,11,-4),
		to_sfixed(3.84,11,-4),
		to_sfixed(2.12,11,-4),
		to_sfixed(18.8,11,-4),
		to_sfixed(90,11,-4),
		to_sfixed(2.45,11,-4),
		to_sfixed(2.68,11,-4),
		to_sfixed(0.27,11,-4),
		to_sfixed(1.48,11,-4),
		to_sfixed(4.28,11,-4),
		to_sfixed(0.91,11,-4),
		to_sfixed(3,11,-4),
		to_sfixed(1035,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.88,11,-4),
		to_sfixed(1.89,11,-4),
		to_sfixed(2.59,11,-4),
		to_sfixed(15,11,-4),
		to_sfixed(101,11,-4),
		to_sfixed(3.25,11,-4),
		to_sfixed(3.56,11,-4),
		to_sfixed(0.17,11,-4),
		to_sfixed(1.7,11,-4),
		to_sfixed(5.43,11,-4),
		to_sfixed(0.88,11,-4),
		to_sfixed(3.56,11,-4),
		to_sfixed(1095,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.24,11,-4),
		to_sfixed(3.98,11,-4),
		to_sfixed(2.29,11,-4),
		to_sfixed(17.5,11,-4),
		to_sfixed(103,11,-4),
		to_sfixed(2.64,11,-4),
		to_sfixed(2.63,11,-4),
		to_sfixed(0.32,11,-4),
		to_sfixed(1.66,11,-4),
		to_sfixed(4.36,11,-4),
		to_sfixed(0.82,11,-4),
		to_sfixed(3,11,-4),
		to_sfixed(680,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.05,11,-4),
		to_sfixed(1.77,11,-4),
		to_sfixed(2.10,11,-4),
		to_sfixed(17,11,-4),
		to_sfixed(107,11,-4),
		to_sfixed(3,11,-4),
		to_sfixed(3,11,-4),
		to_sfixed(0.28,11,-4),
		to_sfixed(2.03,11,-4),
		to_sfixed(5.04,11,-4),
		to_sfixed(0.88,11,-4),
		to_sfixed(3.35,11,-4),
		to_sfixed(885,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(14.21,11,-4),
		to_sfixed(4.04,11,-4),
		to_sfixed(2.44,11,-4),
		to_sfixed(18.9,11,-4),
		to_sfixed(111,11,-4),
		to_sfixed(2.85,11,-4),
		to_sfixed(2.65,11,-4),
		to_sfixed(0.3,11,-4),
		to_sfixed(1.25,11,-4),
		to_sfixed(5.24,11,-4),
		to_sfixed(0.87,11,-4),
		to_sfixed(3.33,11,-4),
		to_sfixed(1080,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(14.38,11,-4),
		to_sfixed(3.59,11,-4),
		to_sfixed(2.28,11,-4),
		to_sfixed(16,11,-4),
		to_sfixed(102,11,-4),
		to_sfixed(3.25,11,-4),
		to_sfixed(3.17,11,-4),
		to_sfixed(0.27,11,-4),
		to_sfixed(2.19,11,-4),
		to_sfixed(4.9,11,-4),
		to_sfixed(1.04,11,-4),
		to_sfixed(3.44,11,-4),
		to_sfixed(1065,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.9,11,-4),
		to_sfixed(1.68,11,-4),
		to_sfixed(2.12,11,-4),
		to_sfixed(16,11,-4),
		to_sfixed(101,11,-4),
		to_sfixed(3.1,11,-4),
		to_sfixed(3.39,11,-4),
		to_sfixed(0.21,11,-4),
		to_sfixed(2.14,11,-4),
		to_sfixed(6.1,11,-4),
		to_sfixed(0.91,11,-4),
		to_sfixed(3.33,11,-4),
		to_sfixed(985,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(14.1,11,-4),
		to_sfixed(2.02,11,-4),
		to_sfixed(2.40,11,-4),
		to_sfixed(18.8,11,-4),
		to_sfixed(103,11,-4),
		to_sfixed(2.75,11,-4),
		to_sfixed(2.92,11,-4),
		to_sfixed(0.32,11,-4),
		to_sfixed(2.38,11,-4),
		to_sfixed(6.2,11,-4),
		to_sfixed(1.07,11,-4),
		to_sfixed(2.75,11,-4),
		to_sfixed(1060,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.94,11,-4),
		to_sfixed(1.73,11,-4),
		to_sfixed(2.27,11,-4),
		to_sfixed(17.4,11,-4),
		to_sfixed(108,11,-4),
		to_sfixed(2.88,11,-4),
		to_sfixed(3.54,11,-4),
		to_sfixed(0.32,11,-4),
		to_sfixed(2.08,11,-4),
		to_sfixed(8.90,11,-4),
		to_sfixed(1.12,11,-4),
		to_sfixed(3.1,11,-4),
		to_sfixed(1260,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.05,11,-4),
		to_sfixed(1.73,11,-4),
		to_sfixed(2.04,11,-4),
		to_sfixed(12.4,11,-4),
		to_sfixed(92,11,-4),
		to_sfixed(2.72,11,-4),
		to_sfixed(3.27,11,-4),
		to_sfixed(0.17,11,-4),
		to_sfixed(2.91,11,-4),
		to_sfixed(7.2,11,-4),
		to_sfixed(1.12,11,-4),
		to_sfixed(2.91,11,-4),
		to_sfixed(1150,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.83,11,-4),
		to_sfixed(1.65,11,-4),
		to_sfixed(2.60,11,-4),
		to_sfixed(17.2,11,-4),
		to_sfixed(94,11,-4),
		to_sfixed(2.45,11,-4),
		to_sfixed(2.99,11,-4),
		to_sfixed(0.22,11,-4),
		to_sfixed(2.29,11,-4),
		to_sfixed(5.6,11,-4),
		to_sfixed(1.24,11,-4),
		to_sfixed(3.37,11,-4),
		to_sfixed(1265,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.82,11,-4),
		to_sfixed(1.75,11,-4),
		to_sfixed(2.42,11,-4),
		to_sfixed(14,11,-4),
		to_sfixed(111,11,-4),
		to_sfixed(3.88,11,-4),
		to_sfixed(3.74,11,-4),
		to_sfixed(0.32,11,-4),
		to_sfixed(1.87,11,-4),
		to_sfixed(7.05,11,-4),
		to_sfixed(1.01,11,-4),
		to_sfixed(3.26,11,-4),
		to_sfixed(1190,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.77,11,-4),
		to_sfixed(1.90,11,-4),
		to_sfixed(2.68,11,-4),
		to_sfixed(17.1,11,-4),
		to_sfixed(115,11,-4),
		to_sfixed(3,11,-4),
		to_sfixed(2.79,11,-4),
		to_sfixed(0.39,11,-4),
		to_sfixed(1.68,11,-4),
		to_sfixed(6.3,11,-4),
		to_sfixed(1.13,11,-4),
		to_sfixed(2.93,11,-4),
		to_sfixed(1375,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.74,11,-4),
		to_sfixed(1.67,11,-4),
		to_sfixed(2.25,11,-4),
		to_sfixed(16.4,11,-4),
		to_sfixed(118,11,-4),
		to_sfixed(2.6,11,-4),
		to_sfixed(2.9,11,-4),
		to_sfixed(0.21,11,-4),
		to_sfixed(1.62,11,-4),
		to_sfixed(5.85,11,-4),
		to_sfixed(0.92,11,-4),
		to_sfixed(3.2,11,-4),
		to_sfixed(1060,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.56,11,-4),
		to_sfixed(1.73,11,-4),
		to_sfixed(2.46,11,-4),
		to_sfixed(20.5,11,-4),
		to_sfixed(116,11,-4),
		to_sfixed(2.96,11,-4),
		to_sfixed(2.78,11,-4),
		to_sfixed(0.2,11,-4),
		to_sfixed(2.45,11,-4),
		to_sfixed(6.25,11,-4),
		to_sfixed(0.98,11,-4),
		to_sfixed(3.03,11,-4),
		to_sfixed(1120,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(14.22,11,-4),
		to_sfixed(1.70,11,-4),
		to_sfixed(2.30,11,-4),
		to_sfixed(16.3,11,-4),
		to_sfixed(118,11,-4),
		to_sfixed(3.2,11,-4),
		to_sfixed(3,11,-4),
		to_sfixed(0.26,11,-4),
		to_sfixed(2.03,11,-4),
		to_sfixed(6.38,11,-4),
		to_sfixed(0.94,11,-4),
		to_sfixed(3.31,11,-4),
		to_sfixed(970,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.29,11,-4),
		to_sfixed(1.97,11,-4),
		to_sfixed(2.68,11,-4),
		to_sfixed(16.8,11,-4),
		to_sfixed(102,11,-4),
		to_sfixed(3,11,-4),
		to_sfixed(3.23,11,-4),
		to_sfixed(0.31,11,-4),
		to_sfixed(1.66,11,-4),
		to_sfixed(6,11,-4),
		to_sfixed(1.07,11,-4),
		to_sfixed(2.84,11,-4),
		to_sfixed(1270,11,-4)
		),

		(
		to_sfixed(1,11,-4),
		to_sfixed(13.72,11,-4),
		to_sfixed(1.43,11,-4),
		to_sfixed(2.50,11,-4),
		to_sfixed(16.7,11,-4),
		to_sfixed(108,11,-4),
		to_sfixed(3.4,11,-4),
		to_sfixed(3.67,11,-4),
		to_sfixed(0.19,11,-4),
		to_sfixed(2.04,11,-4),
		to_sfixed(6.8,11,-4),
		to_sfixed(0.89,11,-4),
		to_sfixed(2.87,11,-4),
		to_sfixed(1285,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.37,11,-4),
		to_sfixed(0.94,11,-4),
		to_sfixed(1.36,11,-4),
		to_sfixed(10.6,11,-4),
		to_sfixed(88,11,-4),
		to_sfixed(1.98,11,-4),
		to_sfixed(0.57,11,-4),
		to_sfixed(0.28,11,-4),
		to_sfixed(0.42,11,-4),
		to_sfixed(1.95,11,-4),
		to_sfixed(1.05,11,-4),
		to_sfixed(1.82,11,-4),
		to_sfixed(520,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.33,11,-4),
		to_sfixed(1.10,11,-4),
		to_sfixed(2.28,11,-4),
		to_sfixed(16,11,-4),
		to_sfixed(101,11,-4),
		to_sfixed(2.05,11,-4),
		to_sfixed(1.09,11,-4),
		to_sfixed(0.63,11,-4),
		to_sfixed(0.41,11,-4),
		to_sfixed(3.27,11,-4),
		to_sfixed(1.25,11,-4),
		to_sfixed(1.67,11,-4),
		to_sfixed(680,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.64,11,-4),
		to_sfixed(1.36,11,-4),
		to_sfixed(2.02,11,-4),
		to_sfixed(16.8,11,-4),
		to_sfixed(100,11,-4),
		to_sfixed(2.02,11,-4),
		to_sfixed(1.41,11,-4),
		to_sfixed(0.53,11,-4),
		to_sfixed(0.62,11,-4),
		to_sfixed(5.75,11,-4),
		to_sfixed(0.98,11,-4),
		to_sfixed(1.59,11,-4),
		to_sfixed(450,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(13.67,11,-4),
		to_sfixed(1.25,11,-4),
		to_sfixed(1.92,11,-4),
		to_sfixed(18,11,-4),
		to_sfixed(94,11,-4),
		to_sfixed(2.1,11,-4),
		to_sfixed(1.79,11,-4),
		to_sfixed(0.32,11,-4),
		to_sfixed(0.73,11,-4),
		to_sfixed(3.8,11,-4),
		to_sfixed(1.23,11,-4),
		to_sfixed(2.46,11,-4),
		to_sfixed(630,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.37,11,-4),
		to_sfixed(1.13,11,-4),
		to_sfixed(2.16,11,-4),
		to_sfixed(19,11,-4),
		to_sfixed(87,11,-4),
		to_sfixed(3.5,11,-4),
		to_sfixed(3.1,11,-4),
		to_sfixed(0.19,11,-4),
		to_sfixed(1.87,11,-4),
		to_sfixed(4.45,11,-4),
		to_sfixed(1.22,11,-4),
		to_sfixed(2.87,11,-4),
		to_sfixed(420,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.17,11,-4),
		to_sfixed(1.45,11,-4),
		to_sfixed(2.53,11,-4),
		to_sfixed(19,11,-4),
		to_sfixed(104,11,-4),
		to_sfixed(1.89,11,-4),
		to_sfixed(1.75,11,-4),
		to_sfixed(0.45,11,-4),
		to_sfixed(1.03,11,-4),
		to_sfixed(2.95,11,-4),
		to_sfixed(1.45,11,-4),
		to_sfixed(2.23,11,-4),
		to_sfixed(355,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.37,11,-4),
		to_sfixed(1.21,11,-4),
		to_sfixed(2.56,11,-4),
		to_sfixed(18.1,11,-4),
		to_sfixed(98,11,-4),
		to_sfixed(2.42,11,-4),
		to_sfixed(2.65,11,-4),
		to_sfixed(0.37,11,-4),
		to_sfixed(2.08,11,-4),
		to_sfixed(4.6,11,-4),
		to_sfixed(1.19,11,-4),
		to_sfixed(2.3,11,-4),
		to_sfixed(678,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(13.11,11,-4),
		to_sfixed(1.01,11,-4),
		to_sfixed(1.70,11,-4),
		to_sfixed(15,11,-4),
		to_sfixed(78,11,-4),
		to_sfixed(2.98,11,-4),
		to_sfixed(3.18,11,-4),
		to_sfixed(0.26,11,-4),
		to_sfixed(2.28,11,-4),
		to_sfixed(5.3,11,-4),
		to_sfixed(1.12,11,-4),
		to_sfixed(3.18,11,-4),
		to_sfixed(502,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.37,11,-4),
		to_sfixed(1.17,11,-4),
		to_sfixed(1.92,11,-4),
		to_sfixed(19.6,11,-4),
		to_sfixed(78,11,-4),
		to_sfixed(2.11,11,-4),
		to_sfixed(2,11,-4),
		to_sfixed(0.27,11,-4),
		to_sfixed(1.04,11,-4),
		to_sfixed(4.68,11,-4),
		to_sfixed(1.12,11,-4),
		to_sfixed(3.48,11,-4),
		to_sfixed(510,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(13.34,11,-4),
		to_sfixed(0.94,11,-4),
		to_sfixed(2.36,11,-4),
		to_sfixed(17,11,-4),
		to_sfixed(110,11,-4),
		to_sfixed(2.53,11,-4),
		to_sfixed(1.3,11,-4),
		to_sfixed(0.55,11,-4),
		to_sfixed(0.42,11,-4),
		to_sfixed(3.17,11,-4),
		to_sfixed(1.02,11,-4),
		to_sfixed(1.93,11,-4),
		to_sfixed(750,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.21,11,-4),
		to_sfixed(1.19,11,-4),
		to_sfixed(1.75,11,-4),
		to_sfixed(16.8,11,-4),
		to_sfixed(151,11,-4),
		to_sfixed(1.85,11,-4),
		to_sfixed(1.28,11,-4),
		to_sfixed(0.14,11,-4),
		to_sfixed(2.5,11,-4),
		to_sfixed(2.85,11,-4),
		to_sfixed(1.28,11,-4),
		to_sfixed(3.07,11,-4),
		to_sfixed(718,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.29,11,-4),
		to_sfixed(1.61,11,-4),
		to_sfixed(2.21,11,-4),
		to_sfixed(20.4,11,-4),
		to_sfixed(103,11,-4),
		to_sfixed(1.1,11,-4),
		to_sfixed(1.02,11,-4),
		to_sfixed(0.37,11,-4),
		to_sfixed(1.46,11,-4),
		to_sfixed(3.05,11,-4),
		to_sfixed(0.906,11,-4),
		to_sfixed(1.82,11,-4),
		to_sfixed(870,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(13.86,11,-4),
		to_sfixed(1.51,11,-4),
		to_sfixed(2.67,11,-4),
		to_sfixed(25,11,-4),
		to_sfixed(86,11,-4),
		to_sfixed(2.95,11,-4),
		to_sfixed(2.86,11,-4),
		to_sfixed(0.21,11,-4),
		to_sfixed(1.87,11,-4),
		to_sfixed(3.38,11,-4),
		to_sfixed(1.36,11,-4),
		to_sfixed(3.16,11,-4),
		to_sfixed(410,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(13.49,11,-4),
		to_sfixed(1.66,11,-4),
		to_sfixed(2.24,11,-4),
		to_sfixed(24,11,-4),
		to_sfixed(87,11,-4),
		to_sfixed(1.88,11,-4),
		to_sfixed(1.84,11,-4),
		to_sfixed(0.27,11,-4),
		to_sfixed(1.03,11,-4),
		to_sfixed(3.74,11,-4),
		to_sfixed(0.98,11,-4),
		to_sfixed(2.78,11,-4),
		to_sfixed(472,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.99,11,-4),
		to_sfixed(1.67,11,-4),
		to_sfixed(2.60,11,-4),
		to_sfixed(30,11,-4),
		to_sfixed(139,11,-4),
		to_sfixed(3.3,11,-4),
		to_sfixed(2.89,11,-4),
		to_sfixed(0.21,11,-4),
		to_sfixed(1.96,11,-4),
		to_sfixed(3.35,11,-4),
		to_sfixed(1.31,11,-4),
		to_sfixed(3.5,11,-4),
		to_sfixed(985,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(11.96,11,-4),
		to_sfixed(1.09,11,-4),
		to_sfixed(2.30,11,-4),
		to_sfixed(21,11,-4),
		to_sfixed(101,11,-4),
		to_sfixed(3.38,11,-4),
		to_sfixed(2.14,11,-4),
		to_sfixed(0.13,11,-4),
		to_sfixed(1.65,11,-4),
		to_sfixed(3.21,11,-4),
		to_sfixed(0.99,11,-4),
		to_sfixed(3.13,11,-4),
		to_sfixed(886,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(11.66,11,-4),
		to_sfixed(1.88,11,-4),
		to_sfixed(1.92,11,-4),
		to_sfixed(16,11,-4),
		to_sfixed(97,11,-4),
		to_sfixed(1.61,11,-4),
		to_sfixed(1.57,11,-4),
		to_sfixed(0.34,11,-4),
		to_sfixed(1.15,11,-4),
		to_sfixed(3.8,11,-4),
		to_sfixed(1.23,11,-4),
		to_sfixed(2.14,11,-4),
		to_sfixed(428,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(13.03,11,-4),
		to_sfixed(0.90,11,-4),
		to_sfixed(1.71,11,-4),
		to_sfixed(16,11,-4),
		to_sfixed(86,11,-4),
		to_sfixed(1.95,11,-4),
		to_sfixed(2.03,11,-4),
		to_sfixed(0.24,11,-4),
		to_sfixed(1.46,11,-4),
		to_sfixed(4.6,11,-4),
		to_sfixed(1.19,11,-4),
		to_sfixed(2.48,11,-4),
		to_sfixed(392,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(11.84,11,-4),
		to_sfixed(2.89,11,-4),
		to_sfixed(2.23,11,-4),
		to_sfixed(18,11,-4),
		to_sfixed(112,11,-4),
		to_sfixed(1.72,11,-4),
		to_sfixed(1.32,11,-4),
		to_sfixed(0.43,11,-4),
		to_sfixed(0.95,11,-4),
		to_sfixed(2.65,11,-4),
		to_sfixed(0.96,11,-4),
		to_sfixed(2.52,11,-4),
		to_sfixed(500,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.33,11,-4),
		to_sfixed(0.99,11,-4),
		to_sfixed(1.95,11,-4),
		to_sfixed(14.8,11,-4),
		to_sfixed(136,11,-4),
		to_sfixed(1.9,11,-4),
		to_sfixed(1.85,11,-4),
		to_sfixed(0.35,11,-4),
		to_sfixed(2.76,11,-4),
		to_sfixed(3.4,11,-4),
		to_sfixed(1.06,11,-4),
		to_sfixed(2.31,11,-4),
		to_sfixed(750,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.7,11,-4),
		to_sfixed(3.87,11,-4),
		to_sfixed(2.40,11,-4),
		to_sfixed(23,11,-4),
		to_sfixed(101,11,-4),
		to_sfixed(2.83,11,-4),
		to_sfixed(2.55,11,-4),
		to_sfixed(0.43,11,-4),
		to_sfixed(1.95,11,-4),
		to_sfixed(2.57,11,-4),
		to_sfixed(1.19,11,-4),
		to_sfixed(3.13,11,-4),
		to_sfixed(463,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12,11,-4),
		to_sfixed(0.92,11,-4),
		to_sfixed(2,11,-4),
		to_sfixed(19,11,-4),
		to_sfixed(86,11,-4),
		to_sfixed(2.42,11,-4),
		to_sfixed(2.26,11,-4),
		to_sfixed(0.3,11,-4),
		to_sfixed(1.43,11,-4),
		to_sfixed(2.5,11,-4),
		to_sfixed(1.38,11,-4),
		to_sfixed(3.12,11,-4),
		to_sfixed(278,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.72,11,-4),
		to_sfixed(1.81,11,-4),
		to_sfixed(2.20,11,-4),
		to_sfixed(18.8,11,-4),
		to_sfixed(86,11,-4),
		to_sfixed(2.2,11,-4),
		to_sfixed(2.53,11,-4),
		to_sfixed(0.26,11,-4),
		to_sfixed(1.77,11,-4),
		to_sfixed(3.9,11,-4),
		to_sfixed(1.16,11,-4),
		to_sfixed(3.14,11,-4),
		to_sfixed(714,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.08,11,-4),
		to_sfixed(1.13,11,-4),
		to_sfixed(2.51,11,-4),
		to_sfixed(24,11,-4),
		to_sfixed(78,11,-4),
		to_sfixed(2,11,-4),
		to_sfixed(1.58,11,-4),
		to_sfixed(0.4,11,-4),
		to_sfixed(1.4,11,-4),
		to_sfixed(2.2,11,-4),
		to_sfixed(1.31,11,-4),
		to_sfixed(2.72,11,-4),
		to_sfixed(630,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(13.05,11,-4),
		to_sfixed(3.86,11,-4),
		to_sfixed(2.32,11,-4),
		to_sfixed(22.5,11,-4),
		to_sfixed(85,11,-4),
		to_sfixed(1.65,11,-4),
		to_sfixed(1.59,11,-4),
		to_sfixed(0.61,11,-4),
		to_sfixed(1.62,11,-4),
		to_sfixed(4.8,11,-4),
		to_sfixed(0.84,11,-4),
		to_sfixed(2.01,11,-4),
		to_sfixed(515,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(11.84,11,-4),
		to_sfixed(0.89,11,-4),
		to_sfixed(2.58,11,-4),
		to_sfixed(18,11,-4),
		to_sfixed(94,11,-4),
		to_sfixed(2.2,11,-4),
		to_sfixed(2.21,11,-4),
		to_sfixed(0.22,11,-4),
		to_sfixed(2.35,11,-4),
		to_sfixed(3.05,11,-4),
		to_sfixed(0.79,11,-4),
		to_sfixed(3.08,11,-4),
		to_sfixed(520,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.67,11,-4),
		to_sfixed(0.98,11,-4),
		to_sfixed(2.24,11,-4),
		to_sfixed(18,11,-4),
		to_sfixed(99,11,-4),
		to_sfixed(2.2,11,-4),
		to_sfixed(1.94,11,-4),
		to_sfixed(0.3,11,-4),
		to_sfixed(1.46,11,-4),
		to_sfixed(2.62,11,-4),
		to_sfixed(1.23,11,-4),
		to_sfixed(3.16,11,-4),
		to_sfixed(450,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.16,11,-4),
		to_sfixed(1.61,11,-4),
		to_sfixed(2.31,11,-4),
		to_sfixed(22.8,11,-4),
		to_sfixed(90,11,-4),
		to_sfixed(1.78,11,-4),
		to_sfixed(1.69,11,-4),
		to_sfixed(0.43,11,-4),
		to_sfixed(1.56,11,-4),
		to_sfixed(2.45,11,-4),
		to_sfixed(1.33,11,-4),
		to_sfixed(2.26,11,-4),
		to_sfixed(495,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(11.65,11,-4),
		to_sfixed(1.67,11,-4),
		to_sfixed(2.62,11,-4),
		to_sfixed(26,11,-4),
		to_sfixed(88,11,-4),
		to_sfixed(1.92,11,-4),
		to_sfixed(1.61,11,-4),
		to_sfixed(0.4,11,-4),
		to_sfixed(1.34,11,-4),
		to_sfixed(2.6,11,-4),
		to_sfixed(1.36,11,-4),
		to_sfixed(3.21,11,-4),
		to_sfixed(562,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(11.64,11,-4),
		to_sfixed(2.06,11,-4),
		to_sfixed(2.46,11,-4),
		to_sfixed(21.6,11,-4),
		to_sfixed(84,11,-4),
		to_sfixed(1.95,11,-4),
		to_sfixed(1.69,11,-4),
		to_sfixed(0.48,11,-4),
		to_sfixed(1.35,11,-4),
		to_sfixed(2.8,11,-4),
		to_sfixed(1,11,-4),
		to_sfixed(2.75,11,-4),
		to_sfixed(680,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.08,11,-4),
		to_sfixed(1.33,11,-4),
		to_sfixed(2.30,11,-4),
		to_sfixed(23.6,11,-4),
		to_sfixed(70,11,-4),
		to_sfixed(2.2,11,-4),
		to_sfixed(1.59,11,-4),
		to_sfixed(0.42,11,-4),
		to_sfixed(1.38,11,-4),
		to_sfixed(1.74,11,-4),
		to_sfixed(1.07,11,-4),
		to_sfixed(3.21,11,-4),
		to_sfixed(625,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.08,11,-4),
		to_sfixed(1.83,11,-4),
		to_sfixed(2.32,11,-4),
		to_sfixed(18.5,11,-4),
		to_sfixed(81,11,-4),
		to_sfixed(1.6,11,-4),
		to_sfixed(1.5,11,-4),
		to_sfixed(0.52,11,-4),
		to_sfixed(1.64,11,-4),
		to_sfixed(2.4,11,-4),
		to_sfixed(1.08,11,-4),
		to_sfixed(2.27,11,-4),
		to_sfixed(480,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12,11,-4),
		to_sfixed(1.51,11,-4),
		to_sfixed(2.42,11,-4),
		to_sfixed(22,11,-4),
		to_sfixed(86,11,-4),
		to_sfixed(1.45,11,-4),
		to_sfixed(1.25,11,-4),
		to_sfixed(0.5,11,-4),
		to_sfixed(1.63,11,-4),
		to_sfixed(3.6,11,-4),
		to_sfixed(1.05,11,-4),
		to_sfixed(2.65,11,-4),
		to_sfixed(450,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.69,11,-4),
		to_sfixed(1.53,11,-4),
		to_sfixed(2.26,11,-4),
		to_sfixed(20.7,11,-4),
		to_sfixed(80,11,-4),
		to_sfixed(1.38,11,-4),
		to_sfixed(1.46,11,-4),
		to_sfixed(0.58,11,-4),
		to_sfixed(1.62,11,-4),
		to_sfixed(3.05,11,-4),
		to_sfixed(0.96,11,-4),
		to_sfixed(2.06,11,-4),
		to_sfixed(495,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.29,11,-4),
		to_sfixed(2.83,11,-4),
		to_sfixed(2.22,11,-4),
		to_sfixed(18,11,-4),
		to_sfixed(88,11,-4),
		to_sfixed(2.45,11,-4),
		to_sfixed(2.25,11,-4),
		to_sfixed(0.25,11,-4),
		to_sfixed(1.99,11,-4),
		to_sfixed(2.15,11,-4),
		to_sfixed(1.15,11,-4),
		to_sfixed(3.3,11,-4),
		to_sfixed(290,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(11.62,11,-4),
		to_sfixed(1.99,11,-4),
		to_sfixed(2.28,11,-4),
		to_sfixed(18,11,-4),
		to_sfixed(98,11,-4),
		to_sfixed(3.02,11,-4),
		to_sfixed(2.26,11,-4),
		to_sfixed(0.17,11,-4),
		to_sfixed(1.35,11,-4),
		to_sfixed(3.25,11,-4),
		to_sfixed(1.16,11,-4),
		to_sfixed(2.96,11,-4),
		to_sfixed(345,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.47,11,-4),
		to_sfixed(1.52,11,-4),
		to_sfixed(2.20,11,-4),
		to_sfixed(19,11,-4),
		to_sfixed(162,11,-4),
		to_sfixed(2.5,11,-4),
		to_sfixed(2.27,11,-4),
		to_sfixed(0.32,11,-4),
		to_sfixed(3.28,11,-4),
		to_sfixed(2.6,11,-4),
		to_sfixed(1.16,11,-4),
		to_sfixed(2.63,11,-4),
		to_sfixed(937,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(11.81,11,-4),
		to_sfixed(2.12,11,-4),
		to_sfixed(2.74,11,-4),
		to_sfixed(21.5,11,-4),
		to_sfixed(134,11,-4),
		to_sfixed(1.6,11,-4),
		to_sfixed(0.99,11,-4),
		to_sfixed(0.14,11,-4),
		to_sfixed(1.56,11,-4),
		to_sfixed(2.5,11,-4),
		to_sfixed(0.95,11,-4),
		to_sfixed(2.26,11,-4),
		to_sfixed(625,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.29,11,-4),
		to_sfixed(1.41,11,-4),
		to_sfixed(1.98,11,-4),
		to_sfixed(16,11,-4),
		to_sfixed(85,11,-4),
		to_sfixed(2.55,11,-4),
		to_sfixed(2.5,11,-4),
		to_sfixed(0.29,11,-4),
		to_sfixed(1.77,11,-4),
		to_sfixed(2.9,11,-4),
		to_sfixed(1.23,11,-4),
		to_sfixed(2.74,11,-4),
		to_sfixed(428,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.37,11,-4),
		to_sfixed(1.07,11,-4),
		to_sfixed(2.10,11,-4),
		to_sfixed(18.5,11,-4),
		to_sfixed(88,11,-4),
		to_sfixed(3.52,11,-4),
		to_sfixed(3.75,11,-4),
		to_sfixed(0.24,11,-4),
		to_sfixed(1.95,11,-4),
		to_sfixed(4.5,11,-4),
		to_sfixed(1.04,11,-4),
		to_sfixed(2.77,11,-4),
		to_sfixed(660,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.29,11,-4),
		to_sfixed(3.17,11,-4),
		to_sfixed(2.21,11,-4),
		to_sfixed(18,11,-4),
		to_sfixed(88,11,-4),
		to_sfixed(2.85,11,-4),
		to_sfixed(2.99,11,-4),
		to_sfixed(0.45,11,-4),
		to_sfixed(2.81,11,-4),
		to_sfixed(2.3,11,-4),
		to_sfixed(1.42,11,-4),
		to_sfixed(2.83,11,-4),
		to_sfixed(406,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.08,11,-4),
		to_sfixed(2.08,11,-4),
		to_sfixed(1.70,11,-4),
		to_sfixed(17.5,11,-4),
		to_sfixed(97,11,-4),
		to_sfixed(2.23,11,-4),
		to_sfixed(2.17,11,-4),
		to_sfixed(0.26,11,-4),
		to_sfixed(1.4,11,-4),
		to_sfixed(3.3,11,-4),
		to_sfixed(1.27,11,-4),
		to_sfixed(2.96,11,-4),
		to_sfixed(710,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.6,11,-4),
		to_sfixed(1.34,11,-4),
		to_sfixed(1.90,11,-4),
		to_sfixed(18.5,11,-4),
		to_sfixed(88,11,-4),
		to_sfixed(1.45,11,-4),
		to_sfixed(1.36,11,-4),
		to_sfixed(0.29,11,-4),
		to_sfixed(1.35,11,-4),
		to_sfixed(2.45,11,-4),
		to_sfixed(1.04,11,-4),
		to_sfixed(2.77,11,-4),
		to_sfixed(562,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.34,11,-4),
		to_sfixed(2.45,11,-4),
		to_sfixed(2.46,11,-4),
		to_sfixed(21,11,-4),
		to_sfixed(98,11,-4),
		to_sfixed(2.56,11,-4),
		to_sfixed(2.11,11,-4),
		to_sfixed(0.34,11,-4),
		to_sfixed(1.31,11,-4),
		to_sfixed(2.8,11,-4),
		to_sfixed(0.8,11,-4),
		to_sfixed(3.38,11,-4),
		to_sfixed(438,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(11.82,11,-4),
		to_sfixed(1.72,11,-4),
		to_sfixed(1.88,11,-4),
		to_sfixed(19.5,11,-4),
		to_sfixed(86,11,-4),
		to_sfixed(2.5,11,-4),
		to_sfixed(1.64,11,-4),
		to_sfixed(0.37,11,-4),
		to_sfixed(1.42,11,-4),
		to_sfixed(2.06,11,-4),
		to_sfixed(0.94,11,-4),
		to_sfixed(2.44,11,-4),
		to_sfixed(415,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.51,11,-4),
		to_sfixed(1.73,11,-4),
		to_sfixed(1.98,11,-4),
		to_sfixed(20.5,11,-4),
		to_sfixed(85,11,-4),
		to_sfixed(2.2,11,-4),
		to_sfixed(1.92,11,-4),
		to_sfixed(0.32,11,-4),
		to_sfixed(1.48,11,-4),
		to_sfixed(2.94,11,-4),
		to_sfixed(1.04,11,-4),
		to_sfixed(3.57,11,-4),
		to_sfixed(672,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.42,11,-4),
		to_sfixed(2.55,11,-4),
		to_sfixed(2.27,11,-4),
		to_sfixed(22,11,-4),
		to_sfixed(90,11,-4),
		to_sfixed(1.68,11,-4),
		to_sfixed(1.84,11,-4),
		to_sfixed(0.66,11,-4),
		to_sfixed(1.42,11,-4),
		to_sfixed(2.7,11,-4),
		to_sfixed(0.86,11,-4),
		to_sfixed(3.3,11,-4),
		to_sfixed(315,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.25,11,-4),
		to_sfixed(1.73,11,-4),
		to_sfixed(2.12,11,-4),
		to_sfixed(19,11,-4),
		to_sfixed(80,11,-4),
		to_sfixed(1.65,11,-4),
		to_sfixed(2.03,11,-4),
		to_sfixed(0.37,11,-4),
		to_sfixed(1.63,11,-4),
		to_sfixed(3.4,11,-4),
		to_sfixed(1,11,-4),
		to_sfixed(3.17,11,-4),
		to_sfixed(510,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.72,11,-4),
		to_sfixed(1.75,11,-4),
		to_sfixed(2.28,11,-4),
		to_sfixed(22.5,11,-4),
		to_sfixed(84,11,-4),
		to_sfixed(1.38,11,-4),
		to_sfixed(1.76,11,-4),
		to_sfixed(0.48,11,-4),
		to_sfixed(1.63,11,-4),
		to_sfixed(3.3,11,-4),
		to_sfixed(0.88,11,-4),
		to_sfixed(2.42,11,-4),
		to_sfixed(488,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.22,11,-4),
		to_sfixed(1.29,11,-4),
		to_sfixed(1.94,11,-4),
		to_sfixed(19,11,-4),
		to_sfixed(92,11,-4),
		to_sfixed(2.36,11,-4),
		to_sfixed(2.04,11,-4),
		to_sfixed(0.39,11,-4),
		to_sfixed(2.08,11,-4),
		to_sfixed(2.7,11,-4),
		to_sfixed(0.86,11,-4),
		to_sfixed(3.02,11,-4),
		to_sfixed(312,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(11.61,11,-4),
		to_sfixed(1.35,11,-4),
		to_sfixed(2.70,11,-4),
		to_sfixed(20,11,-4),
		to_sfixed(94,11,-4),
		to_sfixed(2.74,11,-4),
		to_sfixed(2.92,11,-4),
		to_sfixed(0.29,11,-4),
		to_sfixed(2.49,11,-4),
		to_sfixed(2.65,11,-4),
		to_sfixed(0.96,11,-4),
		to_sfixed(3.26,11,-4),
		to_sfixed(680,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(11.46,11,-4),
		to_sfixed(3.74,11,-4),
		to_sfixed(1.82,11,-4),
		to_sfixed(19.5,11,-4),
		to_sfixed(107,11,-4),
		to_sfixed(3.18,11,-4),
		to_sfixed(2.58,11,-4),
		to_sfixed(0.24,11,-4),
		to_sfixed(3.58,11,-4),
		to_sfixed(2.9,11,-4),
		to_sfixed(0.75,11,-4),
		to_sfixed(2.81,11,-4),
		to_sfixed(562,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.52,11,-4),
		to_sfixed(2.43,11,-4),
		to_sfixed(2.17,11,-4),
		to_sfixed(21,11,-4),
		to_sfixed(88,11,-4),
		to_sfixed(2.55,11,-4),
		to_sfixed(2.27,11,-4),
		to_sfixed(0.26,11,-4),
		to_sfixed(1.22,11,-4),
		to_sfixed(2,11,-4),
		to_sfixed(0.9,11,-4),
		to_sfixed(2.78,11,-4),
		to_sfixed(325,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(11.76,11,-4),
		to_sfixed(2.68,11,-4),
		to_sfixed(2.92,11,-4),
		to_sfixed(20,11,-4),
		to_sfixed(103,11,-4),
		to_sfixed(1.75,11,-4),
		to_sfixed(2.03,11,-4),
		to_sfixed(0.6,11,-4),
		to_sfixed(1.05,11,-4),
		to_sfixed(3.8,11,-4),
		to_sfixed(1.23,11,-4),
		to_sfixed(2.5,11,-4),
		to_sfixed(607,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(11.41,11,-4),
		to_sfixed(0.74,11,-4),
		to_sfixed(2.50,11,-4),
		to_sfixed(21,11,-4),
		to_sfixed(88,11,-4),
		to_sfixed(2.48,11,-4),
		to_sfixed(2.01,11,-4),
		to_sfixed(0.42,11,-4),
		to_sfixed(1.44,11,-4),
		to_sfixed(3.08,11,-4),
		to_sfixed(1.1,11,-4),
		to_sfixed(2.31,11,-4),
		to_sfixed(434,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.08,11,-4),
		to_sfixed(1.39,11,-4),
		to_sfixed(2.50,11,-4),
		to_sfixed(22.5,11,-4),
		to_sfixed(84,11,-4),
		to_sfixed(2.56,11,-4),
		to_sfixed(2.29,11,-4),
		to_sfixed(0.43,11,-4),
		to_sfixed(1.04,11,-4),
		to_sfixed(2.9,11,-4),
		to_sfixed(0.93,11,-4),
		to_sfixed(3.19,11,-4),
		to_sfixed(385,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(11.03,11,-4),
		to_sfixed(1.51,11,-4),
		to_sfixed(2.20,11,-4),
		to_sfixed(21.5,11,-4),
		to_sfixed(85,11,-4),
		to_sfixed(2.46,11,-4),
		to_sfixed(2.17,11,-4),
		to_sfixed(0.52,11,-4),
		to_sfixed(2.01,11,-4),
		to_sfixed(1.9,11,-4),
		to_sfixed(1.71,11,-4),
		to_sfixed(2.87,11,-4),
		to_sfixed(407,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(11.82,11,-4),
		to_sfixed(1.47,11,-4),
		to_sfixed(1.99,11,-4),
		to_sfixed(20.8,11,-4),
		to_sfixed(86,11,-4),
		to_sfixed(1.98,11,-4),
		to_sfixed(1.6,11,-4),
		to_sfixed(0.3,11,-4),
		to_sfixed(1.53,11,-4),
		to_sfixed(1.95,11,-4),
		to_sfixed(0.95,11,-4),
		to_sfixed(3.33,11,-4),
		to_sfixed(495,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.42,11,-4),
		to_sfixed(1.61,11,-4),
		to_sfixed(2.19,11,-4),
		to_sfixed(22.5,11,-4),
		to_sfixed(108,11,-4),
		to_sfixed(2,11,-4),
		to_sfixed(2.09,11,-4),
		to_sfixed(0.34,11,-4),
		to_sfixed(1.61,11,-4),
		to_sfixed(2.06,11,-4),
		to_sfixed(1.06,11,-4),
		to_sfixed(2.96,11,-4),
		to_sfixed(345,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.77,11,-4),
		to_sfixed(3.43,11,-4),
		to_sfixed(1.98,11,-4),
		to_sfixed(16,11,-4),
		to_sfixed(80,11,-4),
		to_sfixed(1.63,11,-4),
		to_sfixed(1.25,11,-4),
		to_sfixed(0.43,11,-4),
		to_sfixed(0.83,11,-4),
		to_sfixed(3.4,11,-4),
		to_sfixed(0.7,11,-4),
		to_sfixed(2.12,11,-4),
		to_sfixed(372,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12,11,-4),
		to_sfixed(3.43,11,-4),
		to_sfixed(2,11,-4),
		to_sfixed(19,11,-4),
		to_sfixed(87,11,-4),
		to_sfixed(2,11,-4),
		to_sfixed(1.64,11,-4),
		to_sfixed(0.37,11,-4),
		to_sfixed(1.87,11,-4),
		to_sfixed(1.28,11,-4),
		to_sfixed(0.93,11,-4),
		to_sfixed(3.05,11,-4),
		to_sfixed(564,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(11.45,11,-4),
		to_sfixed(2.40,11,-4),
		to_sfixed(2.42,11,-4),
		to_sfixed(20,11,-4),
		to_sfixed(96,11,-4),
		to_sfixed(2.9,11,-4),
		to_sfixed(2.79,11,-4),
		to_sfixed(0.32,11,-4),
		to_sfixed(1.83,11,-4),
		to_sfixed(3.25,11,-4),
		to_sfixed(0.8,11,-4),
		to_sfixed(3.39,11,-4),
		to_sfixed(625,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(11.56,11,-4),
		to_sfixed(2.05,11,-4),
		to_sfixed(3.23,11,-4),
		to_sfixed(28.5,11,-4),
		to_sfixed(119,11,-4),
		to_sfixed(3.18,11,-4),
		to_sfixed(5.08,11,-4),
		to_sfixed(0.47,11,-4),
		to_sfixed(1.87,11,-4),
		to_sfixed(6,11,-4),
		to_sfixed(0.93,11,-4),
		to_sfixed(3.69,11,-4),
		to_sfixed(465,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.42,11,-4),
		to_sfixed(4.43,11,-4),
		to_sfixed(2.73,11,-4),
		to_sfixed(26.5,11,-4),
		to_sfixed(102,11,-4),
		to_sfixed(2.2,11,-4),
		to_sfixed(2.13,11,-4),
		to_sfixed(0.43,11,-4),
		to_sfixed(1.71,11,-4),
		to_sfixed(2.08,11,-4),
		to_sfixed(0.92,11,-4),
		to_sfixed(3.12,11,-4),
		to_sfixed(365,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(13.05,11,-4),
		to_sfixed(5.80,11,-4),
		to_sfixed(2.13,11,-4),
		to_sfixed(21.5,11,-4),
		to_sfixed(86,11,-4),
		to_sfixed(2.62,11,-4),
		to_sfixed(2.65,11,-4),
		to_sfixed(0.3,11,-4),
		to_sfixed(2.01,11,-4),
		to_sfixed(2.6,11,-4),
		to_sfixed(0.73,11,-4),
		to_sfixed(3.1,11,-4),
		to_sfixed(380,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(11.87,11,-4),
		to_sfixed(4.31,11,-4),
		to_sfixed(2.39,11,-4),
		to_sfixed(21,11,-4),
		to_sfixed(82,11,-4),
		to_sfixed(2.86,11,-4),
		to_sfixed(3.03,11,-4),
		to_sfixed(0.21,11,-4),
		to_sfixed(2.91,11,-4),
		to_sfixed(2.8,11,-4),
		to_sfixed(0.75,11,-4),
		to_sfixed(3.64,11,-4),
		to_sfixed(380,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.07,11,-4),
		to_sfixed(2.16,11,-4),
		to_sfixed(2.17,11,-4),
		to_sfixed(21,11,-4),
		to_sfixed(85,11,-4),
		to_sfixed(2.6,11,-4),
		to_sfixed(2.65,11,-4),
		to_sfixed(0.37,11,-4),
		to_sfixed(1.35,11,-4),
		to_sfixed(2.76,11,-4),
		to_sfixed(0.86,11,-4),
		to_sfixed(3.28,11,-4),
		to_sfixed(378,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.43,11,-4),
		to_sfixed(1.53,11,-4),
		to_sfixed(2.29,11,-4),
		to_sfixed(21.5,11,-4),
		to_sfixed(86,11,-4),
		to_sfixed(2.74,11,-4),
		to_sfixed(3.15,11,-4),
		to_sfixed(0.39,11,-4),
		to_sfixed(1.77,11,-4),
		to_sfixed(3.94,11,-4),
		to_sfixed(0.69,11,-4),
		to_sfixed(2.84,11,-4),
		to_sfixed(352,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(11.79,11,-4),
		to_sfixed(2.13,11,-4),
		to_sfixed(2.78,11,-4),
		to_sfixed(28.5,11,-4),
		to_sfixed(92,11,-4),
		to_sfixed(2.13,11,-4),
		to_sfixed(2.24,11,-4),
		to_sfixed(0.58,11,-4),
		to_sfixed(1.76,11,-4),
		to_sfixed(3,11,-4),
		to_sfixed(0.97,11,-4),
		to_sfixed(2.44,11,-4),
		to_sfixed(466,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.37,11,-4),
		to_sfixed(1.63,11,-4),
		to_sfixed(2.30,11,-4),
		to_sfixed(24.5,11,-4),
		to_sfixed(88,11,-4),
		to_sfixed(2.22,11,-4),
		to_sfixed(2.45,11,-4),
		to_sfixed(0.4,11,-4),
		to_sfixed(1.9,11,-4),
		to_sfixed(2.12,11,-4),
		to_sfixed(0.89,11,-4),
		to_sfixed(2.78,11,-4),
		to_sfixed(342,11,-4)
		),

		(
		to_sfixed(2,11,-4),
		to_sfixed(12.04,11,-4),
		to_sfixed(4.30,11,-4),
		to_sfixed(2.38,11,-4),
		to_sfixed(22,11,-4),
		to_sfixed(80,11,-4),
		to_sfixed(2.1,11,-4),
		to_sfixed(1.75,11,-4),
		to_sfixed(0.42,11,-4),
		to_sfixed(1.35,11,-4),
		to_sfixed(2.6,11,-4),
		to_sfixed(0.79,11,-4),
		to_sfixed(2.57,11,-4),
		to_sfixed(580,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.86,11,-4),
		to_sfixed(1.35,11,-4),
		to_sfixed(2.32,11,-4),
		to_sfixed(18,11,-4),
		to_sfixed(122,11,-4),
		to_sfixed(1.51,11,-4),
		to_sfixed(1.25,11,-4),
		to_sfixed(0.21,11,-4),
		to_sfixed(0.94,11,-4),
		to_sfixed(4.1,11,-4),
		to_sfixed(0.76,11,-4),
		to_sfixed(1.29,11,-4),
		to_sfixed(630,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.88,11,-4),
		to_sfixed(2.99,11,-4),
		to_sfixed(2.40,11,-4),
		to_sfixed(20,11,-4),
		to_sfixed(104,11,-4),
		to_sfixed(1.3,11,-4),
		to_sfixed(1.22,11,-4),
		to_sfixed(0.24,11,-4),
		to_sfixed(0.83,11,-4),
		to_sfixed(5.4,11,-4),
		to_sfixed(0.74,11,-4),
		to_sfixed(1.42,11,-4),
		to_sfixed(530,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.81,11,-4),
		to_sfixed(2.31,11,-4),
		to_sfixed(2.40,11,-4),
		to_sfixed(24,11,-4),
		to_sfixed(98,11,-4),
		to_sfixed(1.15,11,-4),
		to_sfixed(1.09,11,-4),
		to_sfixed(0.27,11,-4),
		to_sfixed(0.83,11,-4),
		to_sfixed(5.7,11,-4),
		to_sfixed(0.66,11,-4),
		to_sfixed(1.36,11,-4),
		to_sfixed(560,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.7,11,-4),
		to_sfixed(3.55,11,-4),
		to_sfixed(2.36,11,-4),
		to_sfixed(21.5,11,-4),
		to_sfixed(106,11,-4),
		to_sfixed(1.7,11,-4),
		to_sfixed(1.2,11,-4),
		to_sfixed(0.17,11,-4),
		to_sfixed(0.84,11,-4),
		to_sfixed(5,11,-4),
		to_sfixed(0.78,11,-4),
		to_sfixed(1.29,11,-4),
		to_sfixed(600,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.51,11,-4),
		to_sfixed(1.24,11,-4),
		to_sfixed(2.25,11,-4),
		to_sfixed(17.5,11,-4),
		to_sfixed(85,11,-4),
		to_sfixed(2,11,-4),
		to_sfixed(0.58,11,-4),
		to_sfixed(0.6,11,-4),
		to_sfixed(1.25,11,-4),
		to_sfixed(5.45,11,-4),
		to_sfixed(0.75,11,-4),
		to_sfixed(1.51,11,-4),
		to_sfixed(650,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.6,11,-4),
		to_sfixed(2.46,11,-4),
		to_sfixed(2.20,11,-4),
		to_sfixed(18.5,11,-4),
		to_sfixed(94,11,-4),
		to_sfixed(1.62,11,-4),
		to_sfixed(0.66,11,-4),
		to_sfixed(0.63,11,-4),
		to_sfixed(0.94,11,-4),
		to_sfixed(7.1,11,-4),
		to_sfixed(0.73,11,-4),
		to_sfixed(1.58,11,-4),
		to_sfixed(695,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.25,11,-4),
		to_sfixed(4.72,11,-4),
		to_sfixed(2.54,11,-4),
		to_sfixed(21,11,-4),
		to_sfixed(89,11,-4),
		to_sfixed(1.38,11,-4),
		to_sfixed(0.47,11,-4),
		to_sfixed(0.53,11,-4),
		to_sfixed(0.8,11,-4),
		to_sfixed(3.85,11,-4),
		to_sfixed(0.75,11,-4),
		to_sfixed(1.27,11,-4),
		to_sfixed(720,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.53,11,-4),
		to_sfixed(5.51,11,-4),
		to_sfixed(2.64,11,-4),
		to_sfixed(25,11,-4),
		to_sfixed(96,11,-4),
		to_sfixed(1.79,11,-4),
		to_sfixed(0.6,11,-4),
		to_sfixed(0.63,11,-4),
		to_sfixed(1.1,11,-4),
		to_sfixed(5,11,-4),
		to_sfixed(0.82,11,-4),
		to_sfixed(1.69,11,-4),
		to_sfixed(515,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.49,11,-4),
		to_sfixed(3.59,11,-4),
		to_sfixed(2.19,11,-4),
		to_sfixed(19.5,11,-4),
		to_sfixed(88,11,-4),
		to_sfixed(1.62,11,-4),
		to_sfixed(0.48,11,-4),
		to_sfixed(0.58,11,-4),
		to_sfixed(0.88,11,-4),
		to_sfixed(5.7,11,-4),
		to_sfixed(0.81,11,-4),
		to_sfixed(1.82,11,-4),
		to_sfixed(580,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.84,11,-4),
		to_sfixed(2.96,11,-4),
		to_sfixed(2.61,11,-4),
		to_sfixed(24,11,-4),
		to_sfixed(101,11,-4),
		to_sfixed(2.32,11,-4),
		to_sfixed(0.6,11,-4),
		to_sfixed(0.53,11,-4),
		to_sfixed(0.81,11,-4),
		to_sfixed(4.92,11,-4),
		to_sfixed(0.89,11,-4),
		to_sfixed(2.15,11,-4),
		to_sfixed(590,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.93,11,-4),
		to_sfixed(2.81,11,-4),
		to_sfixed(2.70,11,-4),
		to_sfixed(21,11,-4),
		to_sfixed(96,11,-4),
		to_sfixed(1.54,11,-4),
		to_sfixed(0.5,11,-4),
		to_sfixed(0.53,11,-4),
		to_sfixed(0.75,11,-4),
		to_sfixed(4.6,11,-4),
		to_sfixed(0.77,11,-4),
		to_sfixed(2.31,11,-4),
		to_sfixed(600,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.36,11,-4),
		to_sfixed(2.56,11,-4),
		to_sfixed(2.35,11,-4),
		to_sfixed(20,11,-4),
		to_sfixed(89,11,-4),
		to_sfixed(1.4,11,-4),
		to_sfixed(0.5,11,-4),
		to_sfixed(0.37,11,-4),
		to_sfixed(0.64,11,-4),
		to_sfixed(5.6,11,-4),
		to_sfixed(0.7,11,-4),
		to_sfixed(2.47,11,-4),
		to_sfixed(780,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.52,11,-4),
		to_sfixed(3.17,11,-4),
		to_sfixed(2.72,11,-4),
		to_sfixed(23.5,11,-4),
		to_sfixed(97,11,-4),
		to_sfixed(1.55,11,-4),
		to_sfixed(0.52,11,-4),
		to_sfixed(0.5,11,-4),
		to_sfixed(0.55,11,-4),
		to_sfixed(4.35,11,-4),
		to_sfixed(0.89,11,-4),
		to_sfixed(2.06,11,-4),
		to_sfixed(520,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.62,11,-4),
		to_sfixed(4.95,11,-4),
		to_sfixed(2.35,11,-4),
		to_sfixed(20,11,-4),
		to_sfixed(92,11,-4),
		to_sfixed(2,11,-4),
		to_sfixed(0.8,11,-4),
		to_sfixed(0.47,11,-4),
		to_sfixed(1.02,11,-4),
		to_sfixed(4.4,11,-4),
		to_sfixed(0.91,11,-4),
		to_sfixed(2.05,11,-4),
		to_sfixed(550,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.25,11,-4),
		to_sfixed(3.88,11,-4),
		to_sfixed(2.20,11,-4),
		to_sfixed(18.5,11,-4),
		to_sfixed(112,11,-4),
		to_sfixed(1.38,11,-4),
		to_sfixed(0.78,11,-4),
		to_sfixed(0.29,11,-4),
		to_sfixed(1.14,11,-4),
		to_sfixed(8.21,11,-4),
		to_sfixed(0.65,11,-4),
		to_sfixed(2,11,-4),
		to_sfixed(855,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.16,11,-4),
		to_sfixed(3.57,11,-4),
		to_sfixed(2.15,11,-4),
		to_sfixed(21,11,-4),
		to_sfixed(102,11,-4),
		to_sfixed(1.5,11,-4),
		to_sfixed(0.55,11,-4),
		to_sfixed(0.43,11,-4),
		to_sfixed(1.3,11,-4),
		to_sfixed(4,11,-4),
		to_sfixed(0.6,11,-4),
		to_sfixed(1.68,11,-4),
		to_sfixed(830,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.88,11,-4),
		to_sfixed(5.04,11,-4),
		to_sfixed(2.23,11,-4),
		to_sfixed(20,11,-4),
		to_sfixed(80,11,-4),
		to_sfixed(0.98,11,-4),
		to_sfixed(0.34,11,-4),
		to_sfixed(0.4,11,-4),
		to_sfixed(0.68,11,-4),
		to_sfixed(4.9,11,-4),
		to_sfixed(0.58,11,-4),
		to_sfixed(1.33,11,-4),
		to_sfixed(415,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.87,11,-4),
		to_sfixed(4.61,11,-4),
		to_sfixed(2.48,11,-4),
		to_sfixed(21.5,11,-4),
		to_sfixed(86,11,-4),
		to_sfixed(1.7,11,-4),
		to_sfixed(0.65,11,-4),
		to_sfixed(0.47,11,-4),
		to_sfixed(0.86,11,-4),
		to_sfixed(7.65,11,-4),
		to_sfixed(0.54,11,-4),
		to_sfixed(1.86,11,-4),
		to_sfixed(625,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.32,11,-4),
		to_sfixed(3.24,11,-4),
		to_sfixed(2.38,11,-4),
		to_sfixed(21.5,11,-4),
		to_sfixed(92,11,-4),
		to_sfixed(1.93,11,-4),
		to_sfixed(0.76,11,-4),
		to_sfixed(0.45,11,-4),
		to_sfixed(1.25,11,-4),
		to_sfixed(8.42,11,-4),
		to_sfixed(0.55,11,-4),
		to_sfixed(1.62,11,-4),
		to_sfixed(650,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.08,11,-4),
		to_sfixed(3.90,11,-4),
		to_sfixed(2.36,11,-4),
		to_sfixed(21.5,11,-4),
		to_sfixed(113,11,-4),
		to_sfixed(1.41,11,-4),
		to_sfixed(1.39,11,-4),
		to_sfixed(0.34,11,-4),
		to_sfixed(1.14,11,-4),
		to_sfixed(9.40,11,-4),
		to_sfixed(0.57,11,-4),
		to_sfixed(1.33,11,-4),
		to_sfixed(550,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.5,11,-4),
		to_sfixed(3.12,11,-4),
		to_sfixed(2.62,11,-4),
		to_sfixed(24,11,-4),
		to_sfixed(123,11,-4),
		to_sfixed(1.4,11,-4),
		to_sfixed(1.57,11,-4),
		to_sfixed(0.22,11,-4),
		to_sfixed(1.25,11,-4),
		to_sfixed(8.60,11,-4),
		to_sfixed(0.59,11,-4),
		to_sfixed(1.3,11,-4),
		to_sfixed(500,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.79,11,-4),
		to_sfixed(2.67,11,-4),
		to_sfixed(2.48,11,-4),
		to_sfixed(22,11,-4),
		to_sfixed(112,11,-4),
		to_sfixed(1.48,11,-4),
		to_sfixed(1.36,11,-4),
		to_sfixed(0.24,11,-4),
		to_sfixed(1.26,11,-4),
		to_sfixed(10.8,11,-4),
		to_sfixed(0.48,11,-4),
		to_sfixed(1.47,11,-4),
		to_sfixed(480,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.11,11,-4),
		to_sfixed(1.90,11,-4),
		to_sfixed(2.75,11,-4),
		to_sfixed(25.5,11,-4),
		to_sfixed(116,11,-4),
		to_sfixed(2.2,11,-4),
		to_sfixed(1.28,11,-4),
		to_sfixed(0.26,11,-4),
		to_sfixed(1.56,11,-4),
		to_sfixed(7.1,11,-4),
		to_sfixed(0.61,11,-4),
		to_sfixed(1.33,11,-4),
		to_sfixed(425,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.23,11,-4),
		to_sfixed(3.30,11,-4),
		to_sfixed(2.28,11,-4),
		to_sfixed(18.5,11,-4),
		to_sfixed(98,11,-4),
		to_sfixed(1.8,11,-4),
		to_sfixed(0.83,11,-4),
		to_sfixed(0.61,11,-4),
		to_sfixed(1.87,11,-4),
		to_sfixed(10.52,11,-4),
		to_sfixed(0.56,11,-4),
		to_sfixed(1.51,11,-4),
		to_sfixed(675,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.58,11,-4),
		to_sfixed(1.29,11,-4),
		to_sfixed(2.10,11,-4),
		to_sfixed(20,11,-4),
		to_sfixed(103,11,-4),
		to_sfixed(1.48,11,-4),
		to_sfixed(0.58,11,-4),
		to_sfixed(0.53,11,-4),
		to_sfixed(1.4,11,-4),
		to_sfixed(7.6,11,-4),
		to_sfixed(0.58,11,-4),
		to_sfixed(1.55,11,-4),
		to_sfixed(640,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.17,11,-4),
		to_sfixed(5.19,11,-4),
		to_sfixed(2.32,11,-4),
		to_sfixed(22,11,-4),
		to_sfixed(93,11,-4),
		to_sfixed(1.74,11,-4),
		to_sfixed(0.63,11,-4),
		to_sfixed(0.61,11,-4),
		to_sfixed(1.55,11,-4),
		to_sfixed(7.9,11,-4),
		to_sfixed(0.6,11,-4),
		to_sfixed(1.48,11,-4),
		to_sfixed(725,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.84,11,-4),
		to_sfixed(4.12,11,-4),
		to_sfixed(2.38,11,-4),
		to_sfixed(19.5,11,-4),
		to_sfixed(89,11,-4),
		to_sfixed(1.8,11,-4),
		to_sfixed(0.83,11,-4),
		to_sfixed(0.48,11,-4),
		to_sfixed(1.56,11,-4),
		to_sfixed(9.01,11,-4),
		to_sfixed(0.57,11,-4),
		to_sfixed(1.64,11,-4),
		to_sfixed(480,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.45,11,-4),
		to_sfixed(3.03,11,-4),
		to_sfixed(2.64,11,-4),
		to_sfixed(27,11,-4),
		to_sfixed(97,11,-4),
		to_sfixed(1.9,11,-4),
		to_sfixed(0.58,11,-4),
		to_sfixed(0.63,11,-4),
		to_sfixed(1.14,11,-4),
		to_sfixed(7.5,11,-4),
		to_sfixed(0.67,11,-4),
		to_sfixed(1.73,11,-4),
		to_sfixed(880,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(14.34,11,-4),
		to_sfixed(1.68,11,-4),
		to_sfixed(2.70,11,-4),
		to_sfixed(25,11,-4),
		to_sfixed(98,11,-4),
		to_sfixed(2.8,11,-4),
		to_sfixed(1.31,11,-4),
		to_sfixed(0.53,11,-4),
		to_sfixed(2.7,11,-4),
		to_sfixed(13,11,-4),
		to_sfixed(0.57,11,-4),
		to_sfixed(1.96,11,-4),
		to_sfixed(660,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.48,11,-4),
		to_sfixed(1.67,11,-4),
		to_sfixed(2.64,11,-4),
		to_sfixed(22.5,11,-4),
		to_sfixed(89,11,-4),
		to_sfixed(2.6,11,-4),
		to_sfixed(1.1,11,-4),
		to_sfixed(0.52,11,-4),
		to_sfixed(2.29,11,-4),
		to_sfixed(11.75,11,-4),
		to_sfixed(0.57,11,-4),
		to_sfixed(1.78,11,-4),
		to_sfixed(620,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.36,11,-4),
		to_sfixed(3.83,11,-4),
		to_sfixed(2.38,11,-4),
		to_sfixed(21,11,-4),
		to_sfixed(88,11,-4),
		to_sfixed(2.3,11,-4),
		to_sfixed(0.92,11,-4),
		to_sfixed(0.5,11,-4),
		to_sfixed(1.04,11,-4),
		to_sfixed(7.65,11,-4),
		to_sfixed(0.56,11,-4),
		to_sfixed(1.58,11,-4),
		to_sfixed(520,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.69,11,-4),
		to_sfixed(3.26,11,-4),
		to_sfixed(2.54,11,-4),
		to_sfixed(20,11,-4),
		to_sfixed(107,11,-4),
		to_sfixed(1.83,11,-4),
		to_sfixed(0.56,11,-4),
		to_sfixed(0.5,11,-4),
		to_sfixed(0.8,11,-4),
		to_sfixed(5.88,11,-4),
		to_sfixed(0.96,11,-4),
		to_sfixed(1.82,11,-4),
		to_sfixed(680,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.85,11,-4),
		to_sfixed(3.27,11,-4),
		to_sfixed(2.58,11,-4),
		to_sfixed(22,11,-4),
		to_sfixed(106,11,-4),
		to_sfixed(1.65,11,-4),
		to_sfixed(0.6,11,-4),
		to_sfixed(0.6,11,-4),
		to_sfixed(0.96,11,-4),
		to_sfixed(5.58,11,-4),
		to_sfixed(0.87,11,-4),
		to_sfixed(2.11,11,-4),
		to_sfixed(570,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.96,11,-4),
		to_sfixed(3.45,11,-4),
		to_sfixed(2.35,11,-4),
		to_sfixed(18.5,11,-4),
		to_sfixed(106,11,-4),
		to_sfixed(1.39,11,-4),
		to_sfixed(0.7,11,-4),
		to_sfixed(0.4,11,-4),
		to_sfixed(0.94,11,-4),
		to_sfixed(5.28,11,-4),
		to_sfixed(0.68,11,-4),
		to_sfixed(1.75,11,-4),
		to_sfixed(675,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.78,11,-4),
		to_sfixed(2.76,11,-4),
		to_sfixed(2.30,11,-4),
		to_sfixed(22,11,-4),
		to_sfixed(90,11,-4),
		to_sfixed(1.35,11,-4),
		to_sfixed(0.68,11,-4),
		to_sfixed(0.41,11,-4),
		to_sfixed(1.03,11,-4),
		to_sfixed(9.58,11,-4),
		to_sfixed(0.7,11,-4),
		to_sfixed(1.68,11,-4),
		to_sfixed(615,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.73,11,-4),
		to_sfixed(4.36,11,-4),
		to_sfixed(2.26,11,-4),
		to_sfixed(22.5,11,-4),
		to_sfixed(88,11,-4),
		to_sfixed(1.28,11,-4),
		to_sfixed(0.47,11,-4),
		to_sfixed(0.52,11,-4),
		to_sfixed(1.15,11,-4),
		to_sfixed(6.62,11,-4),
		to_sfixed(0.78,11,-4),
		to_sfixed(1.75,11,-4),
		to_sfixed(520,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.45,11,-4),
		to_sfixed(3.70,11,-4),
		to_sfixed(2.60,11,-4),
		to_sfixed(23,11,-4),
		to_sfixed(111,11,-4),
		to_sfixed(1.7,11,-4),
		to_sfixed(0.92,11,-4),
		to_sfixed(0.43,11,-4),
		to_sfixed(1.46,11,-4),
		to_sfixed(10.68,11,-4),
		to_sfixed(0.85,11,-4),
		to_sfixed(1.56,11,-4),
		to_sfixed(695,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.82,11,-4),
		to_sfixed(3.37,11,-4),
		to_sfixed(2.30,11,-4),
		to_sfixed(19.5,11,-4),
		to_sfixed(88,11,-4),
		to_sfixed(1.48,11,-4),
		to_sfixed(0.66,11,-4),
		to_sfixed(0.4,11,-4),
		to_sfixed(0.97,11,-4),
		to_sfixed(10.26,11,-4),
		to_sfixed(0.72,11,-4),
		to_sfixed(1.75,11,-4),
		to_sfixed(685,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.58,11,-4),
		to_sfixed(2.58,11,-4),
		to_sfixed(2.69,11,-4),
		to_sfixed(24.5,11,-4),
		to_sfixed(105,11,-4),
		to_sfixed(1.55,11,-4),
		to_sfixed(0.84,11,-4),
		to_sfixed(0.39,11,-4),
		to_sfixed(1.54,11,-4),
		to_sfixed(8.66,11,-4),
		to_sfixed(0.74,11,-4),
		to_sfixed(1.8,11,-4),
		to_sfixed(750,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.4,11,-4),
		to_sfixed(4.60,11,-4),
		to_sfixed(2.86,11,-4),
		to_sfixed(25,11,-4),
		to_sfixed(112,11,-4),
		to_sfixed(1.98,11,-4),
		to_sfixed(0.96,11,-4),
		to_sfixed(0.27,11,-4),
		to_sfixed(1.11,11,-4),
		to_sfixed(8.5,11,-4),
		to_sfixed(0.67,11,-4),
		to_sfixed(1.92,11,-4),
		to_sfixed(630,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.2,11,-4),
		to_sfixed(3.03,11,-4),
		to_sfixed(2.32,11,-4),
		to_sfixed(19,11,-4),
		to_sfixed(96,11,-4),
		to_sfixed(1.25,11,-4),
		to_sfixed(0.49,11,-4),
		to_sfixed(0.4,11,-4),
		to_sfixed(0.73,11,-4),
		to_sfixed(5.5,11,-4),
		to_sfixed(0.66,11,-4),
		to_sfixed(1.83,11,-4),
		to_sfixed(510,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(12.77,11,-4),
		to_sfixed(2.39,11,-4),
		to_sfixed(2.28,11,-4),
		to_sfixed(19.5,11,-4),
		to_sfixed(86,11,-4),
		to_sfixed(1.39,11,-4),
		to_sfixed(0.51,11,-4),
		to_sfixed(0.48,11,-4),
		to_sfixed(0.64,11,-4),
		to_sfixed(9.90,11,-4),
		to_sfixed(0.57,11,-4),
		to_sfixed(1.63,11,-4),
		to_sfixed(470,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(14.16,11,-4),
		to_sfixed(2.51,11,-4),
		to_sfixed(2.48,11,-4),
		to_sfixed(20,11,-4),
		to_sfixed(91,11,-4),
		to_sfixed(1.68,11,-4),
		to_sfixed(0.7,11,-4),
		to_sfixed(0.44,11,-4),
		to_sfixed(1.24,11,-4),
		to_sfixed(9.7,11,-4),
		to_sfixed(0.62,11,-4),
		to_sfixed(1.71,11,-4),
		to_sfixed(660,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.71,11,-4),
		to_sfixed(5.65,11,-4),
		to_sfixed(2.45,11,-4),
		to_sfixed(20.5,11,-4),
		to_sfixed(95,11,-4),
		to_sfixed(1.68,11,-4),
		to_sfixed(0.61,11,-4),
		to_sfixed(0.52,11,-4),
		to_sfixed(1.06,11,-4),
		to_sfixed(7.7,11,-4),
		to_sfixed(0.64,11,-4),
		to_sfixed(1.74,11,-4),
		to_sfixed(740,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.4,11,-4),
		to_sfixed(3.91,11,-4),
		to_sfixed(2.48,11,-4),
		to_sfixed(23,11,-4),
		to_sfixed(102,11,-4),
		to_sfixed(1.8,11,-4),
		to_sfixed(0.75,11,-4),
		to_sfixed(0.43,11,-4),
		to_sfixed(1.41,11,-4),
		to_sfixed(7.3,11,-4),
		to_sfixed(0.7,11,-4),
		to_sfixed(1.56,11,-4),
		to_sfixed(750,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.27,11,-4),
		to_sfixed(4.28,11,-4),
		to_sfixed(2.26,11,-4),
		to_sfixed(20,11,-4),
		to_sfixed(120,11,-4),
		to_sfixed(1.59,11,-4),
		to_sfixed(0.69,11,-4),
		to_sfixed(0.43,11,-4),
		to_sfixed(1.35,11,-4),
		to_sfixed(10.2,11,-4),
		to_sfixed(0.59,11,-4),
		to_sfixed(1.56,11,-4),
		to_sfixed(835,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(13.17,11,-4),
		to_sfixed(2.59,11,-4),
		to_sfixed(2.37,11,-4),
		to_sfixed(20,11,-4),
		to_sfixed(120,11,-4),
		to_sfixed(1.65,11,-4),
		to_sfixed(0.68,11,-4),
		to_sfixed(0.53,11,-4),
		to_sfixed(1.46,11,-4),
		to_sfixed(9.3,11,-4),
		to_sfixed(0.6,11,-4),
		to_sfixed(1.62,11,-4),
		to_sfixed(840,11,-4)
		),

		(
		to_sfixed(3,11,-4),
		to_sfixed(14.13,11,-4),
		to_sfixed(4.10,11,-4),
		to_sfixed(2.74,11,-4),
		to_sfixed(24.5,11,-4),
		to_sfixed(96,11,-4),
		to_sfixed(2.05,11,-4),
		to_sfixed(0.76,11,-4),
		to_sfixed(0.56,11,-4),
		to_sfixed(1.35,11,-4),
		to_sfixed(9.2,11,-4),
		to_sfixed(0.61,11,-4),
		to_sfixed(1.6,11,-4),
		to_sfixed(560,11,-4)
		)

	); 


	
end package body;

    
