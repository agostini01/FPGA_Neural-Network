-------------------------------------------------------
-- Design Name : User Pakage
-- File Name   : neural_net_pkg.vhd
-- Function    : Defines function for LFSR
-- Coder       : Agostini, N. & Barbosa, F.
-------------------------------------------------------
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;

	use work.fixed_float_types.all; -- ieee_proposed for VHDL-93 version
	use work.fixed_pkg.all; -- ieee_proposed for compatibility version

package NN_PKG is

			type INT_ARRAY is array (integer range <>) of integer;
			constant INPUT_PERCEPTRONS 	: integer := 4;
			constant HIDDEN_PERCEPTRONS 	: integer := 4;
			constant OUT_PERCEPTRONS 		: integer := 4;
			constant FIX_SIZE 	: sfixed := to_sfixed(6.5 ,5,-2);
			
			type FIX_ARRAY is array (integer range <>) of sfixed;
			type FIX_ARRAY_2D is array (integer range <>) of FIX_ARRAY;
			type FIX_ARRAY_3D is array (integer range <>) of FIX_ARRAY_2D;

			type T_WINE_DATASET is array (0 to 177, 0 to 12) of sfixed;

end;

package body NN_PKG is
	
	-- biases and weights for input layer
	constant wine_dataset_init_input_layer : FIX_ARRAY_2D(0 to 12) := (
	
	-- biases and weights for hidden layer
		(to_sfixed(1,5,4),to_sfixed(0,5,4)),
		(to_sfixed(1,5,4),to_sfixed(0,5,4)),
		(to_sfixed(1,5,4),to_sfixed(0,5,4)),
		(to_sfixed(1,5,4),to_sfixed(0,5,4)),
		(to_sfixed(1,5,4),to_sfixed(0,5,4)),
		(to_sfixed(1,5,4),to_sfixed(0,5,4)),
		(to_sfixed(1,5,4),to_sfixed(0,5,4)),
		(to_sfixed(1,5,4),to_sfixed(0,5,4)),
		(to_sfixed(1,5,4),to_sfixed(0,5,4)),
		(to_sfixed(1,5,4),to_sfixed(0,5,4)),
		(to_sfixed(1,5,4),to_sfixed(0,5,4)),
		(to_sfixed(1,5,4),to_sfixed(0,5,4)),
		(to_sfixed(1,5,4),to_sfixed(0,5,4))
	);

	constant wine_dataset_init_hidden_layer : FIX_ARRAY_2D(0 to 2) := (
	
	-- biases and weights for output layer
		(to_sfixed(-0.2944,5,4),to_sfixed(-0.1762,5,4),to_sfixed(0.0424,5,4),to_sfixed(0.4687,5,4),to_sfixed(-0.5961,5,4),to_sfixed(-0.7336,5,4),to_sfixed(0.0010,5,4),to_sfixed(-0.4148,5,4),to_sfixed(-0.2067,5,4),to_sfixed(0.1213,5,4),to_sfixed(0.1815,5,4),to_sfixed(-0.3707,5,4),to_sfixed(0.1376,5,4),to_sfixed(2.1061,5,4)),
		(to_sfixed(-1.9218,5,4),to_sfixed(-0.8591,5,4),to_sfixed(-2.2805,5,4),to_sfixed(2.3456,5,4),to_sfixed(-0.1239,5,4),to_sfixed(-0.0335,5,4),to_sfixed(-0.6953,5,4),to_sfixed(0.0853,5,4),to_sfixed(-0.0385,5,4),to_sfixed(-0.4995,5,4),to_sfixed(0.6088,5,4),to_sfixed(-1.4969,5,4),to_sfixed(-2.6136,5,4),to_sfixed(-0.4546,5,4)),
		(to_sfixed(-0.3840,5,4),to_sfixed(-0.6723,5,4),to_sfixed(-0.5043,5,4),to_sfixed(-0.3566,5,4),to_sfixed(-0.0082,5,4),to_sfixed(-0.6894,5,4),to_sfixed(2.8733,5,4),to_sfixed(0.7266,5,4),to_sfixed(1.0385,5,4),to_sfixed(-2.8766,5,4),to_sfixed(1.5652,5,4),to_sfixed(1.8564,5,4),to_sfixed(-0.3278,5,4),to_sfixed(1.9498,5,4))
	);

	constant wine_dataset_init_output_layer : FIX_ARRAY_2D(0 to 2) := (
	
	-- biases and weights matrix
		(to_sfixed(-1.9038,5,4),to_sfixed(-4.1782,5,4),to_sfixed(1.3133,5,4),to_sfixed(0.4581,5,4)),
		(to_sfixed(-1.7035,5,4),to_sfixed(4.1581,5,4),to_sfixed(3.9893,5,4),to_sfixed(-2.2319,5,4)),
		(to_sfixed(0.2439,5,4),to_sfixed(0.0295,5,4),to_sfixed(-4.1666,5,4),to_sfixed(-0.3156,5,4))
	);
	
	constant wine_dataset_init_layer_matrix : FIX_ARRAY_3D(0 to 2) := (
	
	-- wine dataset (https://archive.ics.uci.edu/ml/datasets/Wine)
		(wine_dataset_init_input_layer), 
		(wine_dataset_init_hidden_layer), 
		(wine_dataset_init_output_layer)
	);

	constant wine_dataset : T_WINE_DATASET := (
		(to_sfixed(1,5,4),	to_sfixed(14.23,5,4),	to_sfixed(1.71,5,4),	to_sfixed(2.43,5,4),	to_sfixed(15.6,5,4),	to_sfixed(127,5,4),	to_sfixed(2.8,5,4),	to_sfixed(3.06,5,4),	to_sfixed(0.28,5,4),	to_sfixed(2.29,5,4),	to_sfixed(5.64,5,4),	to_sfixed(1.04,5,4),	to_sfixed(3.92,5,4),	to_sfixed(1065,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.2,5,4),		to_sfixed(1.78,5,4),	to_sfixed(2.14,5,4),	to_sfixed(11.2,5,4),	to_sfixed(100,5,4),	to_sfixed(2.65,5,4),	to_sfixed(2.76,5,4),	to_sfixed(0.26,5,4),	to_sfixed(1.28,5,4),	to_sfixed(4.38,5,4),	to_sfixed(1.05,5,4),	to_sfixed(3.4,5,4),	to_sfixed(1050,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.16,5,4),	to_sfixed(2.36,5,4),	to_sfixed(2.67,5,4),	to_sfixed(18.6,5,4),	to_sfixed(101,5,4),	to_sfixed(2.8,5,4),	to_sfixed(3.24,5,4),	to_sfixed(0.3,5,4),	to_sfixed(2.81,5,4),	to_sfixed(5.68,5,4),	to_sfixed(1.03,5,4),	to_sfixed(3.17,5,4),	to_sfixed(1185,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(14.37,5,4),	to_sfixed(1.95,5,4),	to_sfixed(2.5,5,4),	to_sfixed(16.8,5,4),	to_sfixed(113,5,4),	to_sfixed(3.85,5,4),	to_sfixed(3.49,5,4),	to_sfixed(0.24,5,4),	to_sfixed(2.18,5,4),	to_sfixed(7.8,5,4),	to_sfixed(0.86,5,4),	to_sfixed(3.45,5,4),	to_sfixed(1480,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.24,5,4),	to_sfixed(2.59,5,4),	to_sfixed(2.87,5,4),	to_sfixed(21,5,4),	to_sfixed(118,5,4),	to_sfixed(2.8,5,4),	to_sfixed(2.69,5,4),	to_sfixed(0.39,5,4),	to_sfixed(1.82,5,4),	to_sfixed(4.32,5,4),	to_sfixed(1.04,5,4),	to_sfixed(2.93,5,4),	to_sfixed(735,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(14.2,5,4),		to_sfixed(1.76,5,4),	to_sfixed(2.45,5,4),	to_sfixed(15.2,5,4),	to_sfixed(112,5,4),	to_sfixed(3.27,5,4),	to_sfixed(3.39,5,4),	to_sfixed(0.34,5,4),	to_sfixed(1.97,5,4),	to_sfixed(6.75,5,4),	to_sfixed(1.05,5,4),	to_sfixed(2.85,5,4),	to_sfixed(1450,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(14.39,5,4),	to_sfixed(1.87,5,4),	to_sfixed(2.45,5,4),	to_sfixed(14.6,5,4),	to_sfixed(96,5,4),	to_sfixed(2.5,5,4),	to_sfixed(2.52,5,4),	to_sfixed(0.3,5,4),	to_sfixed(1.98,5,4),	to_sfixed(5.25,5,4),	to_sfixed(1.02,5,4),	to_sfixed(3.58,5,4),	to_sfixed(1290,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(14.06,5,4),	to_sfixed(2.15,5,4),	to_sfixed(2.61,5,4),	to_sfixed(17.6,5,4),	to_sfixed(121,5,4),	to_sfixed(2.6,5,4),	to_sfixed(2.51,5,4),	to_sfixed(0.31,5,4),	to_sfixed(1.25,5,4),	to_sfixed(5.05,5,4),	to_sfixed(1.06,5,4),	to_sfixed(3.58,5,4),	to_sfixed(1295,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(14.83,5,4),	to_sfixed(1.64,5,4),	to_sfixed(2.17,5,4),	to_sfixed(14,5,4),	to_sfixed(97,5,4),	to_sfixed(2.8,5,4),	to_sfixed(2.98,5,4),	to_sfixed(0.29,5,4),	to_sfixed(1.98,5,4),	to_sfixed(5.2,5,4),	to_sfixed(1.08,5,4),	to_sfixed(2.85,5,4),	to_sfixed(1045,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.86,5,4),	to_sfixed(1.35,5,4),	to_sfixed(2.27,5,4),	to_sfixed(16,5,4),	to_sfixed(98,5,4),	to_sfixed(2.98,5,4),	to_sfixed(3.15,5,4),	to_sfixed(0.22,5,4),	to_sfixed(1.85,5,4),	to_sfixed(7.22,5,4),	to_sfixed(1.01,5,4),	to_sfixed(3.55,5,4),	to_sfixed(1045,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(14.1,5,4),		to_sfixed(2.16,5,4),	to_sfixed(2.3,5,4),	to_sfixed(18,5,4),	to_sfixed(105,5,4),	to_sfixed(2.95,5,4),	to_sfixed(3.32,5,4),	to_sfixed(0.22,5,4),	to_sfixed(2.38,5,4),	to_sfixed(5.75,5,4),	to_sfixed(1.25,5,4),	to_sfixed(3.17,5,4),	to_sfixed(1510,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(14.12,5,4),	to_sfixed(1.48,5,4),	to_sfixed(2.32,5,4),	to_sfixed(16.8,5,4),	to_sfixed(95,5,4),	to_sfixed(2.2,5,4),	to_sfixed(2.43,5,4),	to_sfixed(0.26,5,4),	to_sfixed(1.57,5,4),	to_sfixed(5,5,4),		to_sfixed(1.17,5,4),	to_sfixed(2.82,5,4),	to_sfixed(1280,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.75,5,4),	to_sfixed(1.73,5,4),	to_sfixed(2.41,5,4),	to_sfixed(16,5,4),	to_sfixed(89,5,4),	to_sfixed(2.6,5,4),	to_sfixed(2.76,5,4),	to_sfixed(0.29,5,4),	to_sfixed(1.81,5,4),	to_sfixed(5.6,5,4),	to_sfixed(1.15,5,4),	to_sfixed(2.9,5,4),	to_sfixed(1320,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(14.75,5,4),	to_sfixed(1.73,5,4),	to_sfixed(2.39,5,4),	to_sfixed(11.4,5,4),	to_sfixed(91,5,4),	to_sfixed(3.1,5,4),	to_sfixed(3.69,5,4),	to_sfixed(0.43,5,4),	to_sfixed(2.81,5,4),	to_sfixed(5.4,5,4),	to_sfixed(1.25,5,4),	to_sfixed(2.73,5,4),	to_sfixed(1150,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(14.38,5,4),	to_sfixed(1.87,5,4),	to_sfixed(2.38,5,4),	to_sfixed(12,5,4),	to_sfixed(102,5,4),	to_sfixed(3.3,5,4),	to_sfixed(3.64,5,4),	to_sfixed(0.29,5,4),	to_sfixed(2.96,5,4),	to_sfixed(7.5,5,4),	to_sfixed(1.2,5,4),	to_sfixed(3,5,4),		to_sfixed(1547,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.63,5,4),	to_sfixed(1.81,5,4),	to_sfixed(2.7,5,4),	to_sfixed(17.2,5,4),	to_sfixed(112,5,4),	to_sfixed(2.85,5,4),	to_sfixed(2.91,5,4),	to_sfixed(0.3,5,4),	to_sfixed(1.46,5,4),	to_sfixed(7.3,5,4),	to_sfixed(1.28,5,4),	to_sfixed(2.88,5,4),	to_sfixed(1310,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(14.3,5,4),		to_sfixed(1.92,5,4),	to_sfixed(2.72,5,4),	to_sfixed(20,5,4),	to_sfixed(120,5,4),	to_sfixed(2.8,5,4),	to_sfixed(3.14,5,4),	to_sfixed(0.33,5,4),	to_sfixed(1.97,5,4),	to_sfixed(6.2,5,4),	to_sfixed(1.07,5,4),	to_sfixed(2.65,5,4),	to_sfixed(1280,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.83,5,4),	to_sfixed(1.57,5,4),	to_sfixed(2.62,5,4),	to_sfixed(20,5,4),	to_sfixed(115,5,4),	to_sfixed(2.95,5,4),	to_sfixed(3.4,5,4),	to_sfixed(0.4,5,4),	to_sfixed(1.72,5,4),	to_sfixed(6.6,5,4),	to_sfixed(1.13,5,4),	to_sfixed(2.57,5,4),	to_sfixed(1130,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(14.19,5,4),	to_sfixed(1.59,5,4),	to_sfixed(2.48,5,4),	to_sfixed(16.5,5,4),	to_sfixed(108,5,4),	to_sfixed(3.3,5,4),	to_sfixed(3.93,5,4),	to_sfixed(0.32,5,4),	to_sfixed(1.86,5,4),	to_sfixed(8.7,5,4),	to_sfixed(1.23,5,4),	to_sfixed(2.82,5,4),	to_sfixed(1680,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.64,5,4),	to_sfixed(3.1,5,4),	to_sfixed(2.56,5,4),	to_sfixed(15.2,5,4),	to_sfixed(116,5,4),	to_sfixed(2.7,5,4),	to_sfixed(3.03,5,4),	to_sfixed(0.17,5,4),	to_sfixed(1.66,5,4),	to_sfixed(5.1,5,4),	to_sfixed(0.96,5,4),	to_sfixed(3.36,5,4),	to_sfixed(845,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(14.06,5,4),	to_sfixed(1.63,5,4),	to_sfixed(2.28,5,4),	to_sfixed(16,5,4),	to_sfixed(126,5,4),	to_sfixed(3,5,4),		to_sfixed(3.17,5,4),	to_sfixed(0.24,5,4),	to_sfixed(2.1,5,4),	to_sfixed(5.65,5,4),	to_sfixed(1.09,5,4),	to_sfixed(3.71,5,4),	to_sfixed(780,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(12.93,5,4),	to_sfixed(3.8,5,4),	to_sfixed(2.65,5,4),	to_sfixed(18.6,5,4),	to_sfixed(102,5,4),	to_sfixed(2.41,5,4),	to_sfixed(2.41,5,4),	to_sfixed(0.25,5,4),	to_sfixed(1.98,5,4),	to_sfixed(4.5,5,4),	to_sfixed(1.03,5,4),	to_sfixed(3.52,5,4),	to_sfixed(770,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.71,5,4),	to_sfixed(1.86,5,4),	to_sfixed(2.36,5,4),	to_sfixed(16.6,5,4),	to_sfixed(101,5,4),	to_sfixed(2.61,5,4),	to_sfixed(2.88,5,4),	to_sfixed(0.27,5,4),	to_sfixed(1.69,5,4),	to_sfixed(3.8,5,4),	to_sfixed(1.11,5,4),	to_sfixed(4,5,4),		to_sfixed(1035,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(12.85,5,4),	to_sfixed(1.6,5,4),	to_sfixed(2.52,5,4),	to_sfixed(17.8,5,4),	to_sfixed(95,5,4),	to_sfixed(2.48,5,4),	to_sfixed(2.37,5,4),	to_sfixed(0.26,5,4),	to_sfixed(1.46,5,4),	to_sfixed(3.93,5,4),	to_sfixed(1.09,5,4),	to_sfixed(3.63,5,4),	to_sfixed(1015,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.5,5,4),		to_sfixed(1.81,5,4),	to_sfixed(2.61,5,4),	to_sfixed(20,5,4),	to_sfixed(96,5,4),	to_sfixed(2.53,5,4),	to_sfixed(2.61,5,4),	to_sfixed(0.28,5,4),	to_sfixed(1.66,5,4),	to_sfixed(3.52,5,4),	to_sfixed(1.12,5,4),	to_sfixed(3.82,5,4),	to_sfixed(845,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.05,5,4),	to_sfixed(2.05,5,4),	to_sfixed(3.22,5,4),	to_sfixed(25,5,4),	to_sfixed(124,5,4),	to_sfixed(2.63,5,4),	to_sfixed(2.68,5,4),	to_sfixed(0.47,5,4),	to_sfixed(1.92,5,4),	to_sfixed(3.58,5,4),	to_sfixed(1.13,5,4),	to_sfixed(3.2,5,4),	to_sfixed(830,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.39,5,4),	to_sfixed(1.77,5,4),	to_sfixed(2.62,5,4),	to_sfixed(16.1,5,4),	to_sfixed(93,5,4),	to_sfixed(2.85,5,4),	to_sfixed(2.94,5,4),	to_sfixed(0.34,5,4),	to_sfixed(1.45,5,4),	to_sfixed(4.8,5,4),	to_sfixed(0.92,5,4),	to_sfixed(3.22,5,4),	to_sfixed(1195,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.3,5,4),		to_sfixed(1.72,5,4),	to_sfixed(2.14,5,4),	to_sfixed(17,5,4),	to_sfixed(94,5,4),	to_sfixed(2.4,5,4),	to_sfixed(2.19,5,4),	to_sfixed(0.27,5,4),	to_sfixed(1.35,5,4),	to_sfixed(3.95,5,4),	to_sfixed(1.02,5,4),	to_sfixed(2.77,5,4),	to_sfixed(1285,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.87,5,4),	to_sfixed(1.9,5,4),	to_sfixed(2.8,5,4),	to_sfixed(19.4,5,4),	to_sfixed(107,5,4),	to_sfixed(2.95,5,4),	to_sfixed(2.97,5,4),	to_sfixed(0.37,5,4),	to_sfixed(1.76,5,4),	to_sfixed(4.5,5,4),	to_sfixed(1.25,5,4),	to_sfixed(3.4,5,4),	to_sfixed(915,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(14.02,5,4),	to_sfixed(1.68,5,4),	to_sfixed(2.21,5,4),	to_sfixed(16,5,4),	to_sfixed(96,5,4),	to_sfixed(2.65,5,4),	to_sfixed(2.33,5,4),	to_sfixed(0.26,5,4),	to_sfixed(1.98,5,4),	to_sfixed(4.7,5,4),	to_sfixed(1.04,5,4),	to_sfixed(3.59,5,4),	to_sfixed(1035,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.73,5,4),	to_sfixed(1.5,5,4),	to_sfixed(2.7,5,4),	to_sfixed(22.5,5,4),	to_sfixed(101,5,4),	to_sfixed(3,5,4),		to_sfixed(3.25,5,4),	to_sfixed(0.29,5,4),	to_sfixed(2.38,5,4),	to_sfixed(5.7,5,4),	to_sfixed(1.19,5,4),	to_sfixed(2.71,5,4),	to_sfixed(1285,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.58,5,4),	to_sfixed(1.66,5,4),	to_sfixed(2.36,5,4),	to_sfixed(19.1,5,4),	to_sfixed(106,5,4),	to_sfixed(2.86,5,4),	to_sfixed(3.19,5,4),	to_sfixed(0.22,5,4),	to_sfixed(1.95,5,4),	to_sfixed(6.9,5,4),	to_sfixed(1.09,5,4),	to_sfixed(2.88,5,4),	to_sfixed(1515,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.68,5,4),	to_sfixed(1.83,5,4),	to_sfixed(2.36,5,4),	to_sfixed(17.2,5,4),	to_sfixed(104,5,4),	to_sfixed(2.42,5,4),	to_sfixed(2.69,5,4),	to_sfixed(0.42,5,4),	to_sfixed(1.97,5,4),	to_sfixed(3.84,5,4),	to_sfixed(1.23,5,4),	to_sfixed(2.87,5,4),	to_sfixed(990,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.76,5,4),	to_sfixed(1.53,5,4),	to_sfixed(2.7,5,4),	to_sfixed(19.5,5,4),	to_sfixed(132,5,4),	to_sfixed(2.95,5,4),	to_sfixed(2.74,5,4),	to_sfixed(0.5,5,4),	to_sfixed(1.35,5,4),	to_sfixed(5.4,5,4),	to_sfixed(1.25,5,4),	to_sfixed(3,5,4),		to_sfixed(1235,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.51,5,4),	to_sfixed(1.8,5,4),	to_sfixed(2.65,5,4),	to_sfixed(19,5,4),	to_sfixed(110,5,4),	to_sfixed(2.35,5,4),	to_sfixed(2.53,5,4),	to_sfixed(0.29,5,4),	to_sfixed(1.54,5,4),	to_sfixed(4.2,5,4),	to_sfixed(1.1,5,4),	to_sfixed(2.87,5,4),	to_sfixed(1095,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.48,5,4),	to_sfixed(1.81,5,4),	to_sfixed(2.41,5,4),	to_sfixed(20.5,5,4),	to_sfixed(100,5,4),	to_sfixed(2.7,5,4),	to_sfixed(2.98,5,4),	to_sfixed(0.26,5,4),	to_sfixed(1.86,5,4),	to_sfixed(5.1,5,4),	to_sfixed(1.04,5,4),	to_sfixed(3.47,5,4),	to_sfixed(920,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.28,5,4),	to_sfixed(1.64,5,4),	to_sfixed(2.84,5,4),	to_sfixed(15.5,5,4),	to_sfixed(110,5,4),	to_sfixed(2.6,5,4),	to_sfixed(2.68,5,4),	to_sfixed(0.34,5,4),	to_sfixed(1.36,5,4),	to_sfixed(4.6,5,4),	to_sfixed(1.09,5,4),	to_sfixed(2.78,5,4),	to_sfixed(880,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.05,5,4),	to_sfixed(1.65,5,4),	to_sfixed(2.55,5,4),	to_sfixed(18,5,4),	to_sfixed(98,5,4),	to_sfixed(2.45,5,4),	to_sfixed(2.43,5,4),	to_sfixed(0.29,5,4),	to_sfixed(1.44,5,4),	to_sfixed(4.25,5,4),	to_sfixed(1.12,5,4),	to_sfixed(2.51,5,4),	to_sfixed(1105,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.07,5,4),	to_sfixed(1.5,5,4),	to_sfixed(2.1,5,4),	to_sfixed(15.5,5,4),	to_sfixed(98,5,4),	to_sfixed(2.4,5,4),	to_sfixed(2.64,5,4),	to_sfixed(0.28,5,4),	to_sfixed(1.37,5,4),	to_sfixed(3.7,5,4),	to_sfixed(1.18,5,4),	to_sfixed(2.69,5,4),	to_sfixed(1020,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(14.22,5,4),	to_sfixed(3.99,5,4),	to_sfixed(2.51,5,4),	to_sfixed(13.2,5,4),	to_sfixed(128,5,4),	to_sfixed(3,5,4),		to_sfixed(3.04,5,4),	to_sfixed(0.2,5,4),	to_sfixed(2.08,5,4),	to_sfixed(5.1,5,4),	to_sfixed(0.89,5,4),	to_sfixed(3.53,5,4),	to_sfixed(760,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.56,5,4),	to_sfixed(1.71,5,4),	to_sfixed(2.31,5,4),	to_sfixed(16.2,5,4),	to_sfixed(117,5,4),	to_sfixed(3.15,5,4),	to_sfixed(3.29,5,4),	to_sfixed(0.34,5,4),	to_sfixed(2.34,5,4),	to_sfixed(6.13,5,4),	to_sfixed(0.95,5,4),	to_sfixed(3.38,5,4),	to_sfixed(795,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.41,5,4),	to_sfixed(3.84,5,4),	to_sfixed(2.12,5,4),	to_sfixed(18.8,5,4),	to_sfixed(90,5,4),	to_sfixed(2.45,5,4),	to_sfixed(2.68,5,4),	to_sfixed(0.27,5,4),	to_sfixed(1.48,5,4),	to_sfixed(4.28,5,4),	to_sfixed(0.91,5,4),	to_sfixed(3,5,4),		to_sfixed(1035,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.88,5,4),	to_sfixed(1.89,5,4),	to_sfixed(2.59,5,4),	to_sfixed(15,5,4),	to_sfixed(101,5,4),	to_sfixed(3.25,5,4),	to_sfixed(3.56,5,4),	to_sfixed(0.17,5,4),	to_sfixed(1.7,5,4),	to_sfixed(5.43,5,4),	to_sfixed(0.88,5,4),	to_sfixed(3.56,5,4),	to_sfixed(1095,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.24,5,4),	to_sfixed(3.98,5,4),	to_sfixed(2.29,5,4),	to_sfixed(17.5,5,4),	to_sfixed(103,5,4),	to_sfixed(2.64,5,4),	to_sfixed(2.63,5,4),	to_sfixed(0.32,5,4),	to_sfixed(1.66,5,4),	to_sfixed(4.36,5,4),	to_sfixed(0.82,5,4),	to_sfixed(3,5,4),		to_sfixed(680,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.05,5,4),	to_sfixed(1.77,5,4),	to_sfixed(2.1,5,4),	to_sfixed(17,5,4),	to_sfixed(107,5,4),	to_sfixed(3,5,4),		to_sfixed(3,5,4),		to_sfixed(0.28,5,4),	to_sfixed(2.03,5,4),	to_sfixed(5.04,5,4),	to_sfixed(0.88,5,4),	to_sfixed(3.35,5,4),	to_sfixed(885,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(14.21,5,4),	to_sfixed(4.04,5,4),	to_sfixed(2.44,5,4),	to_sfixed(18.9,5,4),	to_sfixed(111,5,4),	to_sfixed(2.85,5,4),	to_sfixed(2.65,5,4),	to_sfixed(0.3,5,4),	to_sfixed(1.25,5,4),	to_sfixed(5.24,5,4),	to_sfixed(0.87,5,4),	to_sfixed(3.33,5,4),	to_sfixed(1080,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(14.38,5,4),	to_sfixed(3.59,5,4),	to_sfixed(2.28,5,4),	to_sfixed(16,5,4),	to_sfixed(102,5,4),	to_sfixed(3.25,5,4),	to_sfixed(3.17,5,4),	to_sfixed(0.27,5,4),	to_sfixed(2.19,5,4),	to_sfixed(4.9,5,4),	to_sfixed(1.04,5,4),	to_sfixed(3.44,5,4),	to_sfixed(1065,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.9,5,4),		to_sfixed(1.68,5,4),	to_sfixed(2.12,5,4),	to_sfixed(16,5,4),	to_sfixed(101,5,4),	to_sfixed(3.1,5,4),	to_sfixed(3.39,5,4),	to_sfixed(0.21,5,4),	to_sfixed(2.14,5,4),	to_sfixed(6.1,5,4),	to_sfixed(0.91,5,4),	to_sfixed(3.33,5,4),	to_sfixed(985,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(14.1,5,4),		to_sfixed(2.02,5,4),	to_sfixed(2.4,5,4),	to_sfixed(18.8,5,4),	to_sfixed(103,5,4),	to_sfixed(2.75,5,4),	to_sfixed(2.92,5,4),	to_sfixed(0.32,5,4),	to_sfixed(2.38,5,4),	to_sfixed(6.2,5,4),	to_sfixed(1.07,5,4),	to_sfixed(2.75,5,4),	to_sfixed(1060,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.94,5,4),	to_sfixed(1.73,5,4),	to_sfixed(2.27,5,4),	to_sfixed(17.4,5,4),	to_sfixed(108,5,4),	to_sfixed(2.88,5,4),	to_sfixed(3.54,5,4),	to_sfixed(0.32,5,4),	to_sfixed(2.08,5,4),	to_sfixed(8.90,5,4),	to_sfixed(1.12,5,4),	to_sfixed(3.1,5,4),	to_sfixed(1260,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.05,5,4),	to_sfixed(1.73,5,4),	to_sfixed(2.04,5,4),	to_sfixed(12.4,5,4),	to_sfixed(92,5,4),	to_sfixed(2.72,5,4),	to_sfixed(3.27,5,4),	to_sfixed(0.17,5,4),	to_sfixed(2.91,5,4),	to_sfixed(7.2,5,4),	to_sfixed(1.12,5,4),	to_sfixed(2.91,5,4),	to_sfixed(1150,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.83,5,4),	to_sfixed(1.65,5,4),	to_sfixed(2.6,5,4),	to_sfixed(17.2,5,4),	to_sfixed(94,5,4),	to_sfixed(2.45,5,4),	to_sfixed(2.99,5,4),	to_sfixed(0.22,5,4),	to_sfixed(2.29,5,4),	to_sfixed(5.6,5,4),	to_sfixed(1.24,5,4),	to_sfixed(3.37,5,4),	to_sfixed(1265,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.82,5,4),	to_sfixed(1.75,5,4),	to_sfixed(2.42,5,4),	to_sfixed(14,5,4),	to_sfixed(111,5,4),	to_sfixed(3.88,5,4),	to_sfixed(3.74,5,4),	to_sfixed(0.32,5,4),	to_sfixed(1.87,5,4),	to_sfixed(7.05,5,4),	to_sfixed(1.01,5,4),	to_sfixed(3.26,5,4),	to_sfixed(1190,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.77,5,4),	to_sfixed(1.9,5,4),	to_sfixed(2.68,5,4),	to_sfixed(17.1,5,4),	to_sfixed(115,5,4),	to_sfixed(3,5,4),		to_sfixed(2.79,5,4),	to_sfixed(0.39,5,4),	to_sfixed(1.68,5,4),	to_sfixed(6.3,5,4),	to_sfixed(1.13,5,4),	to_sfixed(2.93,5,4),	to_sfixed(1375,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.74,5,4),	to_sfixed(1.67,5,4),	to_sfixed(2.25,5,4),	to_sfixed(16.4,5,4),	to_sfixed(118,5,4),	to_sfixed(2.6,5,4),	to_sfixed(2.9,5,4),	to_sfixed(0.21,5,4),	to_sfixed(1.62,5,4),	to_sfixed(5.85,5,4),	to_sfixed(0.92,5,4),	to_sfixed(3.2,5,4),	to_sfixed(1060,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.56,5,4),	to_sfixed(1.73,5,4),	to_sfixed(2.46,5,4),	to_sfixed(20.5,5,4),	to_sfixed(116,5,4),	to_sfixed(2.96,5,4),	to_sfixed(2.78,5,4),	to_sfixed(0.2,5,4),	to_sfixed(2.45,5,4),	to_sfixed(6.25,5,4),	to_sfixed(0.98,5,4),	to_sfixed(3.03,5,4),	to_sfixed(1120,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(14.22,5,4),	to_sfixed(1.7,5,4),	to_sfixed(2.3,5,4),	to_sfixed(16.3,5,4),	to_sfixed(118,5,4),	to_sfixed(3.2,5,4),	to_sfixed(3,5,4),		to_sfixed(0.26,5,4),	to_sfixed(2.03,5,4),	to_sfixed(6.38,5,4),	to_sfixed(0.94,5,4),	to_sfixed(3.31,5,4),	to_sfixed(970,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.29,5,4),	to_sfixed(1.97,5,4),	to_sfixed(2.68,5,4),	to_sfixed(16.8,5,4),	to_sfixed(102,5,4),	to_sfixed(3,5,4),		to_sfixed(3.23,5,4),	to_sfixed(0.31,5,4),	to_sfixed(1.66,5,4),	to_sfixed(6,5,4),		to_sfixed(1.07,5,4),	to_sfixed(2.84,5,4),	to_sfixed(1270,5,4)),
		(to_sfixed(1,5,4),	to_sfixed(13.72,5,4),	to_sfixed(1.43,5,4),	to_sfixed(2.5,5,4),	to_sfixed(16.7,5,4),	to_sfixed(108,5,4),	to_sfixed(3.4,5,4),	to_sfixed(3.67,5,4),	to_sfixed(0.19,5,4),	to_sfixed(2.04,5,4),	to_sfixed(6.8,5,4),	to_sfixed(0.89,5,4),	to_sfixed(2.87,5,4),	to_sfixed(1285,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.37,5,4),	to_sfixed(0.94,5,4),	to_sfixed(1.36,5,4),	to_sfixed(10.6,5,4),	to_sfixed(88,5,4),	to_sfixed(1.98,5,4),	to_sfixed(0.57,5,4),	to_sfixed(0.28,5,4),	to_sfixed(0.42,5,4),	to_sfixed(1.95,5,4),	to_sfixed(1.05,5,4),	to_sfixed(1.82,5,4),	to_sfixed(520,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.33,5,4),	to_sfixed(1.1,5,4),	to_sfixed(2.28,5,4),	to_sfixed(16,5,4),	to_sfixed(101,5,4),	to_sfixed(2.05,5,4),	to_sfixed(1.09,5,4),	to_sfixed(0.63,5,4),	to_sfixed(0.41,5,4),	to_sfixed(3.27,5,4),	to_sfixed(1.25,5,4),	to_sfixed(1.67,5,4),	to_sfixed(680,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.64,5,4),	to_sfixed(1.36,5,4),	to_sfixed(2.02,5,4),	to_sfixed(16.8,5,4),	to_sfixed(100,5,4),	to_sfixed(2.02,5,4),	to_sfixed(1.41,5,4),	to_sfixed(0.53,5,4),	to_sfixed(0.62,5,4),	to_sfixed(5.75,5,4),	to_sfixed(0.98,5,4),	to_sfixed(1.59,5,4),	to_sfixed(450,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(13.67,5,4),	to_sfixed(1.25,5,4),	to_sfixed(1.92,5,4),	to_sfixed(18,5,4),	to_sfixed(94,5,4),	to_sfixed(2.1,5,4),	to_sfixed(1.79,5,4),	to_sfixed(0.32,5,4),	to_sfixed(0.73,5,4),	to_sfixed(3.8,5,4),	to_sfixed(1.23,5,4),	to_sfixed(2.46,5,4),	to_sfixed(630,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.37,5,4),	to_sfixed(1.13,5,4),	to_sfixed(2.16,5,4),	to_sfixed(19,5,4),	to_sfixed(87,5,4),	to_sfixed(3.5,5,4),	to_sfixed(3.1,5,4),	to_sfixed(0.19,5,4),	to_sfixed(1.87,5,4),	to_sfixed(4.45,5,4),	to_sfixed(1.22,5,4),	to_sfixed(2.87,5,4),	to_sfixed(420,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.17,5,4),	to_sfixed(1.45,5,4),	to_sfixed(2.53,5,4),	to_sfixed(19,5,4),	to_sfixed(104,5,4),	to_sfixed(1.89,5,4),	to_sfixed(1.75,5,4),	to_sfixed(0.45,5,4),	to_sfixed(1.03,5,4),	to_sfixed(2.95,5,4),	to_sfixed(1.45,5,4),	to_sfixed(2.23,5,4),	to_sfixed(355,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.37,5,4),	to_sfixed(1.21,5,4),	to_sfixed(2.56,5,4),	to_sfixed(18.1,5,4),	to_sfixed(98,5,4),	to_sfixed(2.42,5,4),	to_sfixed(2.65,5,4),	to_sfixed(0.37,5,4),	to_sfixed(2.08,5,4),	to_sfixed(4.6,5,4),	to_sfixed(1.19,5,4),	to_sfixed(2.3,5,4),	to_sfixed(678,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(13.11,5,4),	to_sfixed(1.01,5,4),	to_sfixed(1.7,5,4),	to_sfixed(15,5,4),	to_sfixed(78,5,4),	to_sfixed(2.98,5,4),	to_sfixed(3.18,5,4),	to_sfixed(0.26,5,4),	to_sfixed(2.28,5,4),	to_sfixed(5.3,5,4),	to_sfixed(1.12,5,4),	to_sfixed(3.18,5,4),	to_sfixed(502,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.37,5,4),	to_sfixed(1.17,5,4),	to_sfixed(1.92,5,4),	to_sfixed(19.6,5,4),	to_sfixed(78,5,4),	to_sfixed(2.11,5,4),	to_sfixed(2,5,4),		to_sfixed(0.27,5,4),	to_sfixed(1.04,5,4),	to_sfixed(4.68,5,4),	to_sfixed(1.12,5,4),	to_sfixed(3.48,5,4),	to_sfixed(510,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(13.34,5,4),	to_sfixed(0.94,5,4),	to_sfixed(2.36,5,4),	to_sfixed(17,5,4),	to_sfixed(110,5,4),	to_sfixed(2.53,5,4),	to_sfixed(1.3,5,4),	to_sfixed(0.55,5,4),	to_sfixed(0.42,5,4),	to_sfixed(3.17,5,4),	to_sfixed(1.02,5,4),	to_sfixed(1.93,5,4),	to_sfixed(750,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.21,5,4),	to_sfixed(1.19,5,4),	to_sfixed(1.75,5,4),	to_sfixed(16.8,5,4),	to_sfixed(151,5,4),	to_sfixed(1.85,5,4),	to_sfixed(1.28,5,4),	to_sfixed(0.14,5,4),	to_sfixed(2.5,5,4),	to_sfixed(2.85,5,4),	to_sfixed(1.28,5,4),	to_sfixed(3.07,5,4),	to_sfixed(718,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.29,5,4),	to_sfixed(1.61,5,4),	to_sfixed(2.21,5,4),	to_sfixed(20.4,5,4),	to_sfixed(103,5,4),	to_sfixed(1.1,5,4),	to_sfixed(1.02,5,4),	to_sfixed(0.37,5,4),	to_sfixed(1.46,5,4),	to_sfixed(3.05,5,4),	to_sfixed(0.906,5,4),to_sfixed(1.82,5,4),	to_sfixed(870,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(13.86,5,4),	to_sfixed(1.51,5,4),	to_sfixed(2.67,5,4),	to_sfixed(25,5,4),	to_sfixed(86,5,4),	to_sfixed(2.95,5,4),	to_sfixed(2.86,5,4),	to_sfixed(0.21,5,4),	to_sfixed(1.87,5,4),	to_sfixed(3.38,5,4),	to_sfixed(1.36,5,4),	to_sfixed(3.16,5,4),	to_sfixed(410,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(13.49,5,4),	to_sfixed(1.66,5,4),	to_sfixed(2.24,5,4),	to_sfixed(24,5,4),	to_sfixed(87,5,4),	to_sfixed(1.88,5,4),	to_sfixed(1.84,5,4),	to_sfixed(0.27,5,4),	to_sfixed(1.03,5,4),	to_sfixed(3.74,5,4),	to_sfixed(0.98,5,4),	to_sfixed(2.78,5,4),	to_sfixed(472,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.99,5,4),	to_sfixed(1.67,5,4),	to_sfixed(2.6,5,4),	to_sfixed(30,5,4),	to_sfixed(139,5,4),	to_sfixed(3.3,5,4),	to_sfixed(2.89,5,4),	to_sfixed(0.21,5,4),	to_sfixed(1.96,5,4),	to_sfixed(3.35,5,4),	to_sfixed(1.31,5,4),	to_sfixed(3.5,5,4),	to_sfixed(985,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(11.96,5,4),	to_sfixed(1.09,5,4),	to_sfixed(2.3,5,4),	to_sfixed(21,5,4),	to_sfixed(101,5,4),	to_sfixed(3.38,5,4),	to_sfixed(2.14,5,4),	to_sfixed(0.13,5,4),	to_sfixed(1.65,5,4),	to_sfixed(3.21,5,4),	to_sfixed(0.99,5,4),	to_sfixed(3.13,5,4),	to_sfixed(886,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(11.66,5,4),	to_sfixed(1.88,5,4),	to_sfixed(1.92,5,4),	to_sfixed(16,5,4),	to_sfixed(97,5,4),	to_sfixed(1.61,5,4),	to_sfixed(1.57,5,4),	to_sfixed(0.34,5,4),	to_sfixed(1.15,5,4),	to_sfixed(3.8,5,4),	to_sfixed(1.23,5,4),	to_sfixed(2.14,5,4),	to_sfixed(428,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(13.03,5,4),	to_sfixed(0.9,5,4),	to_sfixed(1.71,5,4),	to_sfixed(16,5,4),	to_sfixed(86,5,4),	to_sfixed(1.95,5,4),	to_sfixed(2.03,5,4),	to_sfixed(0.24,5,4),	to_sfixed(1.46,5,4),	to_sfixed(4.6,5,4),	to_sfixed(1.19,5,4),	to_sfixed(2.48,5,4),	to_sfixed(392,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(11.84,5,4),	to_sfixed(2.89,5,4),	to_sfixed(2.23,5,4),	to_sfixed(18,5,4),	to_sfixed(112,5,4),	to_sfixed(1.72,5,4),	to_sfixed(1.32,5,4),	to_sfixed(0.43,5,4),	to_sfixed(0.95,5,4),	to_sfixed(2.65,5,4),	to_sfixed(0.96,5,4),	to_sfixed(2.52,5,4),	to_sfixed(500,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.33,5,4),	to_sfixed(0.99,5,4),	to_sfixed(1.95,5,4),	to_sfixed(14.8,5,4),	to_sfixed(136,5,4),	to_sfixed(1.9,5,4),	to_sfixed(1.85,5,4),	to_sfixed(0.35,5,4),	to_sfixed(2.76,5,4),	to_sfixed(3.4,5,4),	to_sfixed(1.06,5,4),	to_sfixed(2.31,5,4),	to_sfixed(750,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.7,5,4),		to_sfixed(3.87,5,4),	to_sfixed(2.4,5,4),	to_sfixed(23,5,4),	to_sfixed(101,5,4),	to_sfixed(2.83,5,4),	to_sfixed(2.55,5,4),	to_sfixed(0.43,5,4),	to_sfixed(1.95,5,4),	to_sfixed(2.57,5,4),	to_sfixed(1.19,5,4),	to_sfixed(3.13,5,4),	to_sfixed(463,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12,5,4),		to_sfixed(0.92,5,4),	to_sfixed(2,5,4),		to_sfixed(19,5,4),	to_sfixed(86,5,4),	to_sfixed(2.42,5,4),	to_sfixed(2.26,5,4),	to_sfixed(0.3,5,4),	to_sfixed(1.43,5,4),	to_sfixed(2.5,5,4),	to_sfixed(1.38,5,4),	to_sfixed(3.12,5,4),	to_sfixed(278,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.72,5,4),	to_sfixed(1.81,5,4),	to_sfixed(2.2,5,4),	to_sfixed(18.8,5,4),	to_sfixed(86,5,4),	to_sfixed(2.2,5,4),	to_sfixed(2.53,5,4),	to_sfixed(0.26,5,4),	to_sfixed(1.77,5,4),	to_sfixed(3.9,5,4),	to_sfixed(1.16,5,4),	to_sfixed(3.14,5,4),	to_sfixed(714,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.08,5,4),	to_sfixed(1.13,5,4),	to_sfixed(2.51,5,4),	to_sfixed(24,5,4),	to_sfixed(78,5,4),	to_sfixed(2,5,4),		to_sfixed(1.58,5,4),	to_sfixed(0.4,5,4),	to_sfixed(1.4,5,4),	to_sfixed(2.2,5,4),	to_sfixed(1.31,5,4),	to_sfixed(2.72,5,4),	to_sfixed(630,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(13.05,5,4),	to_sfixed(3.86,5,4),	to_sfixed(2.32,5,4),	to_sfixed(22.5,5,4),	to_sfixed(85,5,4),	to_sfixed(1.65,5,4),	to_sfixed(1.59,5,4),	to_sfixed(0.61,5,4),	to_sfixed(1.62,5,4),	to_sfixed(4.8,5,4),	to_sfixed(0.84,5,4),	to_sfixed(2.01,5,4),	to_sfixed(515,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(11.84,5,4),	to_sfixed(0.89,5,4),	to_sfixed(2.58,5,4),	to_sfixed(18,5,4),	to_sfixed(94,5,4),	to_sfixed(2.2,5,4),	to_sfixed(2.21,5,4),	to_sfixed(0.22,5,4),	to_sfixed(2.35,5,4),	to_sfixed(3.05,5,4),	to_sfixed(0.79,5,4),	to_sfixed(3.08,5,4),	to_sfixed(520,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.67,5,4),	to_sfixed(0.98,5,4),	to_sfixed(2.24,5,4),	to_sfixed(18,5,4),	to_sfixed(99,5,4),	to_sfixed(2.2,5,4),	to_sfixed(1.94,5,4),	to_sfixed(0.3,5,4),	to_sfixed(1.46,5,4),	to_sfixed(2.62,5,4),	to_sfixed(1.23,5,4),	to_sfixed(3.16,5,4),	to_sfixed(450,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.16,5,4),	to_sfixed(1.61,5,4),	to_sfixed(2.31,5,4),	to_sfixed(22.8,5,4),	to_sfixed(90,5,4),	to_sfixed(1.78,5,4),	to_sfixed(1.69,5,4),	to_sfixed(0.43,5,4),	to_sfixed(1.56,5,4),	to_sfixed(2.45,5,4),	to_sfixed(1.33,5,4),	to_sfixed(2.26,5,4),	to_sfixed(495,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(11.65,5,4),	to_sfixed(1.67,5,4),	to_sfixed(2.62,5,4),	to_sfixed(26,5,4),	to_sfixed(88,5,4),	to_sfixed(1.92,5,4),	to_sfixed(1.61,5,4),	to_sfixed(0.4,5,4),	to_sfixed(1.34,5,4),	to_sfixed(2.6,5,4),	to_sfixed(1.36,5,4),	to_sfixed(3.21,5,4),	to_sfixed(562,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(11.64,5,4),	to_sfixed(2.06,5,4),	to_sfixed(2.46,5,4),	to_sfixed(21.6,5,4),	to_sfixed(84,5,4),	to_sfixed(1.95,5,4),	to_sfixed(1.69,5,4),	to_sfixed(0.48,5,4),	to_sfixed(1.35,5,4),	to_sfixed(2.8,5,4),	to_sfixed(1,5,4),		to_sfixed(2.75,5,4),	to_sfixed(680,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.08,5,4),	to_sfixed(1.33,5,4),	to_sfixed(2.3,5,4),	to_sfixed(23.6,5,4),	to_sfixed(70,5,4),	to_sfixed(2.2,5,4),	to_sfixed(1.59,5,4),	to_sfixed(0.42,5,4),	to_sfixed(1.38,5,4),	to_sfixed(1.74,5,4),	to_sfixed(1.07,5,4),	to_sfixed(3.21,5,4),	to_sfixed(625,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.08,5,4),	to_sfixed(1.83,5,4),	to_sfixed(2.32,5,4),	to_sfixed(18.5,5,4),	to_sfixed(81,5,4),	to_sfixed(1.6,5,4),	to_sfixed(1.5,5,4),	to_sfixed(0.52,5,4),	to_sfixed(1.64,5,4),	to_sfixed(2.4,5,4),	to_sfixed(1.08,5,4),	to_sfixed(2.27,5,4),	to_sfixed(480,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12,5,4),		to_sfixed(1.51,5,4),	to_sfixed(2.42,5,4),	to_sfixed(22,5,4),	to_sfixed(86,5,4),	to_sfixed(1.45,5,4),	to_sfixed(1.25,5,4),	to_sfixed(0.5,5,4),	to_sfixed(1.63,5,4),	to_sfixed(3.6,5,4),	to_sfixed(1.05,5,4),	to_sfixed(2.65,5,4),	to_sfixed(450,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.69,5,4),	to_sfixed(1.53,5,4),	to_sfixed(2.26,5,4),	to_sfixed(20.7,5,4),	to_sfixed(80,5,4),	to_sfixed(1.38,5,4),	to_sfixed(1.46,5,4),	to_sfixed(0.58,5,4),	to_sfixed(1.62,5,4),	to_sfixed(3.05,5,4),	to_sfixed(0.96,5,4),	to_sfixed(2.06,5,4),	to_sfixed(495,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.29,5,4),	to_sfixed(2.83,5,4),	to_sfixed(2.22,5,4),	to_sfixed(18,5,4),	to_sfixed(88,5,4),	to_sfixed(2.45,5,4),	to_sfixed(2.25,5,4),	to_sfixed(0.25,5,4),	to_sfixed(1.99,5,4),	to_sfixed(2.15,5,4),	to_sfixed(1.15,5,4),	to_sfixed(3.3,5,4),	to_sfixed(290,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(11.62,5,4),	to_sfixed(1.99,5,4),	to_sfixed(2.28,5,4),	to_sfixed(18,5,4),	to_sfixed(98,5,4),	to_sfixed(3.02,5,4),	to_sfixed(2.26,5,4),	to_sfixed(0.17,5,4),	to_sfixed(1.35,5,4),	to_sfixed(3.25,5,4),	to_sfixed(1.16,5,4),	to_sfixed(2.96,5,4),	to_sfixed(345,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.47,5,4),	to_sfixed(1.52,5,4),	to_sfixed(2.2,5,4),	to_sfixed(19,5,4),	to_sfixed(162,5,4),	to_sfixed(2.5,5,4),	to_sfixed(2.27,5,4),	to_sfixed(0.32,5,4),	to_sfixed(3.28,5,4),	to_sfixed(2.6,5,4),	to_sfixed(1.16,5,4),	to_sfixed(2.63,5,4),	to_sfixed(937,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(11.81,5,4),	to_sfixed(2.12,5,4),	to_sfixed(2.74,5,4),	to_sfixed(21.5,5,4),	to_sfixed(134,5,4),	to_sfixed(1.6,5,4),	to_sfixed(0.99,5,4),	to_sfixed(0.14,5,4),	to_sfixed(1.56,5,4),	to_sfixed(2.5,5,4),	to_sfixed(0.95,5,4),	to_sfixed(2.26,5,4),	to_sfixed(625,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.29,5,4),	to_sfixed(1.41,5,4),	to_sfixed(1.98,5,4),	to_sfixed(16,5,4),	to_sfixed(85,5,4),	to_sfixed(2.55,5,4),	to_sfixed(2.5,5,4),	to_sfixed(0.29,5,4),	to_sfixed(1.77,5,4),	to_sfixed(2.9,5,4),	to_sfixed(1.23,5,4),	to_sfixed(2.74,5,4),	to_sfixed(428,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.37,5,4),	to_sfixed(1.07,5,4),	to_sfixed(2.1,5,4),	to_sfixed(18.5,5,4),	to_sfixed(88,5,4),	to_sfixed(3.52,5,4),	to_sfixed(3.75,5,4),	to_sfixed(0.24,5,4),	to_sfixed(1.95,5,4),	to_sfixed(4.5,5,4),	to_sfixed(1.04,5,4),	to_sfixed(2.77,5,4),	to_sfixed(660,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.29,5,4),	to_sfixed(3.17,5,4),	to_sfixed(2.21,5,4),	to_sfixed(18,5,4),	to_sfixed(88,5,4),	to_sfixed(2.85,5,4),	to_sfixed(2.99,5,4),	to_sfixed(0.45,5,4),	to_sfixed(2.81,5,4),	to_sfixed(2.3,5,4),	to_sfixed(1.42,5,4),	to_sfixed(2.83,5,4),	to_sfixed(406,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.08,5,4),	to_sfixed(2.08,5,4),	to_sfixed(1.7,5,4),	to_sfixed(17.5,5,4),	to_sfixed(97,5,4),	to_sfixed(2.23,5,4),	to_sfixed(2.17,5,4),	to_sfixed(0.26,5,4),	to_sfixed(1.4,5,4),	to_sfixed(3.3,5,4),	to_sfixed(1.27,5,4),	to_sfixed(2.96,5,4),	to_sfixed(710,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.6,5,4),		to_sfixed(1.34,5,4),	to_sfixed(1.9,5,4),	to_sfixed(18.5,5,4),	to_sfixed(88,5,4),	to_sfixed(1.45,5,4),	to_sfixed(1.36,5,4),	to_sfixed(0.29,5,4),	to_sfixed(1.35,5,4),	to_sfixed(2.45,5,4),	to_sfixed(1.04,5,4),	to_sfixed(2.77,5,4),	to_sfixed(562,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.34,5,4),	to_sfixed(2.45,5,4),	to_sfixed(2.46,5,4),	to_sfixed(21,5,4),	to_sfixed(98,5,4),	to_sfixed(2.56,5,4),	to_sfixed(2.11,5,4),	to_sfixed(0.34,5,4),	to_sfixed(1.31,5,4),	to_sfixed(2.8,5,4),	to_sfixed(0.8,5,4),	to_sfixed(3.38,5,4),	to_sfixed(438,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(11.82,5,4),	to_sfixed(1.72,5,4),	to_sfixed(1.88,5,4),	to_sfixed(19.5,5,4),	to_sfixed(86,5,4),	to_sfixed(2.5,5,4),	to_sfixed(1.64,5,4),	to_sfixed(0.37,5,4),	to_sfixed(1.42,5,4),	to_sfixed(2.06,5,4),	to_sfixed(0.94,5,4),	to_sfixed(2.44,5,4),	to_sfixed(415,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.51,5,4),	to_sfixed(1.73,5,4),	to_sfixed(1.98,5,4),	to_sfixed(20.5,5,4),	to_sfixed(85,5,4),	to_sfixed(2.2,5,4),	to_sfixed(1.92,5,4),	to_sfixed(0.32,5,4),	to_sfixed(1.48,5,4),	to_sfixed(2.94,5,4),	to_sfixed(1.04,5,4),	to_sfixed(3.57,5,4),	to_sfixed(672,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.42,5,4),	to_sfixed(2.55,5,4),	to_sfixed(2.27,5,4),	to_sfixed(22,5,4),	to_sfixed(90,5,4),	to_sfixed(1.68,5,4),	to_sfixed(1.84,5,4),	to_sfixed(0.66,5,4),	to_sfixed(1.42,5,4),	to_sfixed(2.7,5,4),	to_sfixed(0.86,5,4),	to_sfixed(3.3,5,4),	to_sfixed(315,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.25,5,4),	to_sfixed(1.73,5,4),	to_sfixed(2.12,5,4),	to_sfixed(19,5,4),	to_sfixed(80,5,4),	to_sfixed(1.65,5,4),	to_sfixed(2.03,5,4),	to_sfixed(0.37,5,4),	to_sfixed(1.63,5,4),	to_sfixed(3.4,5,4),	to_sfixed(1,5,4),	to_sfixed(3.17,5,4),	to_sfixed(510,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.72,5,4),	to_sfixed(1.75,5,4),	to_sfixed(2.28,5,4),	to_sfixed(22.5,5,4),	to_sfixed(84,5,4),	to_sfixed(1.38,5,4),	to_sfixed(1.76,5,4),	to_sfixed(0.48,5,4),	to_sfixed(1.63,5,4),	to_sfixed(3.3,5,4),	to_sfixed(0.88,5,4),	to_sfixed(2.42,5,4),	to_sfixed(488,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.22,5,4),	to_sfixed(1.29,5,4),	to_sfixed(1.94,5,4),	to_sfixed(19,5,4),	to_sfixed(92,5,4),	to_sfixed(2.36,5,4),	to_sfixed(2.04,5,4),	to_sfixed(0.39,5,4),	to_sfixed(2.08,5,4),	to_sfixed(2.7,5,4),	to_sfixed(0.86,5,4),	to_sfixed(3.02,5,4),	to_sfixed(312,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(11.61,5,4),	to_sfixed(1.35,5,4),	to_sfixed(2.7,5,4),	to_sfixed(20,5,4),	to_sfixed(94,5,4),	to_sfixed(2.74,5,4),	to_sfixed(2.92,5,4),	to_sfixed(0.29,5,4),	to_sfixed(2.49,5,4),	to_sfixed(2.65,5,4),	to_sfixed(0.96,5,4),	to_sfixed(3.26,5,4),	to_sfixed(680,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(11.46,5,4),	to_sfixed(3.74,5,4),	to_sfixed(1.82,5,4),	to_sfixed(19.5,5,4),	to_sfixed(107,5,4),	to_sfixed(3.18,5,4),	to_sfixed(2.58,5,4),	to_sfixed(0.24,5,4),	to_sfixed(3.58,5,4),	to_sfixed(2.9,5,4),	to_sfixed(0.75,5,4),	to_sfixed(2.81,5,4),	to_sfixed(562,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.52,5,4),	to_sfixed(2.43,5,4),	to_sfixed(2.17,5,4),	to_sfixed(21,5,4),	to_sfixed(88,5,4),	to_sfixed(2.55,5,4),	to_sfixed(2.27,5,4),	to_sfixed(0.26,5,4),	to_sfixed(1.22,5,4),	to_sfixed(2,5,4),		to_sfixed(0.9,5,4),	to_sfixed(2.78,5,4),	to_sfixed(325,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(11.76,5,4),	to_sfixed(2.68,5,4),	to_sfixed(2.92,5,4),	to_sfixed(20,5,4),	to_sfixed(103,5,4),	to_sfixed(1.75,5,4),	to_sfixed(2.03,5,4),	to_sfixed(0.6,5,4),	to_sfixed(1.05,5,4),	to_sfixed(3.8,5,4),	to_sfixed(1.23,5,4),	to_sfixed(2.5,5,4),	to_sfixed(607,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(11.41,5,4),	to_sfixed(0.74,5,4),	to_sfixed(2.5,5,4),	to_sfixed(21,5,4),	to_sfixed(88,5,4),	to_sfixed(2.48,5,4),	to_sfixed(2.01,5,4),	to_sfixed(0.42,5,4),	to_sfixed(1.44,5,4),	to_sfixed(3.08,5,4),	to_sfixed(1.1,5,4),	to_sfixed(2.31,5,4),	to_sfixed(434,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.08,5,4),	to_sfixed(1.39,5,4),	to_sfixed(2.5,5,4),	to_sfixed(22.5,5,4),	to_sfixed(84,5,4),	to_sfixed(2.56,5,4),	to_sfixed(2.29,5,4),	to_sfixed(0.43,5,4),	to_sfixed(1.04,5,4),	to_sfixed(2.9,5,4),	to_sfixed(0.93,5,4),	to_sfixed(3.19,5,4),	to_sfixed(385,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(11.03,5,4),	to_sfixed(1.51,5,4),	to_sfixed(2.2,5,4),	to_sfixed(21.5,5,4),	to_sfixed(85,5,4),	to_sfixed(2.46,5,4),	to_sfixed(2.17,5,4),	to_sfixed(0.52,5,4),	to_sfixed(2.01,5,4),	to_sfixed(1.9,5,4),	to_sfixed(1.71,5,4),	to_sfixed(2.87,5,4),	to_sfixed(407,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(11.82,5,4),	to_sfixed(1.47,5,4),	to_sfixed(1.99,5,4),	to_sfixed(20.8,5,4),	to_sfixed(86,5,4),	to_sfixed(1.98,5,4),	to_sfixed(1.6,5,4),	to_sfixed(0.3,5,4),	to_sfixed(1.53,5,4),	to_sfixed(1.95,5,4),	to_sfixed(0.95,5,4),	to_sfixed(3.33,5,4),	to_sfixed(495,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.42,5,4),	to_sfixed(1.61,5,4),	to_sfixed(2.19,5,4),	to_sfixed(22.5,5,4),	to_sfixed(108,5,4),	to_sfixed(2,5,4),		to_sfixed(2.09,5,4),	to_sfixed(0.34,5,4),	to_sfixed(1.61,5,4),	to_sfixed(2.06,5,4),	to_sfixed(1.06,5,4),	to_sfixed(2.96,5,4),	to_sfixed(345,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.77,5,4),	to_sfixed(3.43,5,4),	to_sfixed(1.98,5,4),	to_sfixed(16,5,4),	to_sfixed(80,5,4),	to_sfixed(1.63,5,4),	to_sfixed(1.25,5,4),	to_sfixed(0.43,5,4),	to_sfixed(0.83,5,4),	to_sfixed(3.4,5,4),	to_sfixed(0.7,5,4),	to_sfixed(2.12,5,4),	to_sfixed(372,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12,5,4),		to_sfixed(3.43,5,4),	to_sfixed(2,5,4),		to_sfixed(19,5,4),	to_sfixed(87,5,4),	to_sfixed(2,5,4),		to_sfixed(1.64,5,4),	to_sfixed(0.37,5,4),	to_sfixed(1.87,5,4),	to_sfixed(1.28,5,4),	to_sfixed(0.93,5,4),	to_sfixed(3.05,5,4),	to_sfixed(564,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(11.45,5,4),	to_sfixed(2.4,5,4),	to_sfixed(2.42,5,4),	to_sfixed(20,5,4),	to_sfixed(96,5,4),	to_sfixed(2.9,5,4),	to_sfixed(2.79,5,4),	to_sfixed(0.32,5,4),	to_sfixed(1.83,5,4),	to_sfixed(3.25,5,4),	to_sfixed(0.8,5,4),	to_sfixed(3.39,5,4),	to_sfixed(625,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(11.56,5,4),	to_sfixed(2.05,5,4),	to_sfixed(3.23,5,4),	to_sfixed(28.5,5,4),	to_sfixed(119,5,4),	to_sfixed(3.18,5,4),	to_sfixed(5.08,5,4),	to_sfixed(0.47,5,4),	to_sfixed(1.87,5,4),	to_sfixed(6,5,4),		to_sfixed(0.93,5,4),	to_sfixed(3.69,5,4),	to_sfixed(465,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.42,5,4),	to_sfixed(4.43,5,4),	to_sfixed(2.73,5,4),	to_sfixed(26.5,5,4),	to_sfixed(102,5,4),	to_sfixed(2.2,5,4),	to_sfixed(2.13,5,4),	to_sfixed(0.43,5,4),	to_sfixed(1.71,5,4),	to_sfixed(2.08,5,4),	to_sfixed(0.92,5,4),	to_sfixed(3.12,5,4),	to_sfixed(365,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(13.05,5,4),	to_sfixed(5.8,5,4),	to_sfixed(2.13,5,4),	to_sfixed(21.5,5,4),	to_sfixed(86,5,4),	to_sfixed(2.62,5,4),	to_sfixed(2.65,5,4),	to_sfixed(0.3,5,4),	to_sfixed(2.01,5,4),	to_sfixed(2.6,5,4),	to_sfixed(0.73,5,4),	to_sfixed(3.1,5,4),	to_sfixed(380,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(11.87,5,4),	to_sfixed(4.31,5,4),	to_sfixed(2.39,5,4),	to_sfixed(21,5,4),	to_sfixed(82,5,4),	to_sfixed(2.86,5,4),	to_sfixed(3.03,5,4),	to_sfixed(0.21,5,4),	to_sfixed(2.91,5,4),	to_sfixed(2.8,5,4),	to_sfixed(0.75,5,4),	to_sfixed(3.64,5,4),	to_sfixed(380,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.07,5,4),	to_sfixed(2.16,5,4),	to_sfixed(2.17,5,4),	to_sfixed(21,5,4),	to_sfixed(85,5,4),	to_sfixed(2.6,5,4),	to_sfixed(2.65,5,4),	to_sfixed(0.37,5,4),	to_sfixed(1.35,5,4),	to_sfixed(2.76,5,4),	to_sfixed(0.86,5,4),	to_sfixed(3.28,5,4),	to_sfixed(378,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.43,5,4),	to_sfixed(1.53,5,4),	to_sfixed(2.29,5,4),	to_sfixed(21.5,5,4),	to_sfixed(86,5,4),	to_sfixed(2.74,5,4),	to_sfixed(3.15,5,4),	to_sfixed(0.39,5,4),	to_sfixed(1.77,5,4),	to_sfixed(3.94,5,4),	to_sfixed(0.69,5,4),	to_sfixed(2.84,5,4),	to_sfixed(352,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(11.79,5,4),	to_sfixed(2.13,5,4),	to_sfixed(2.78,5,4),	to_sfixed(28.5,5,4),	to_sfixed(92,5,4),	to_sfixed(2.13,5,4),	to_sfixed(2.24,5,4),	to_sfixed(0.58,5,4),	to_sfixed(1.76,5,4),	to_sfixed(3,5,4),		to_sfixed(0.97,5,4),	to_sfixed(2.44,5,4),	to_sfixed(466,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.37,5,4),	to_sfixed(1.63,5,4),	to_sfixed(2.3,5,4),	to_sfixed(24.5,5,4),	to_sfixed(88,5,4),	to_sfixed(2.22,5,4),	to_sfixed(2.45,5,4),	to_sfixed(0.4,5,4),	to_sfixed(1.9,5,4),	to_sfixed(2.12,5,4),	to_sfixed(0.89,5,4),	to_sfixed(2.78,5,4),	to_sfixed(342,5,4)),
		(to_sfixed(2,5,4),	to_sfixed(12.04,5,4),	to_sfixed(4.3,5,4),	to_sfixed(2.38,5,4),	to_sfixed(22,5,4),	to_sfixed(80,5,4),	to_sfixed(2.1,5,4),	to_sfixed(1.75,5,4),	to_sfixed(0.42,5,4),	to_sfixed(1.35,5,4),	to_sfixed(2.6,5,4),	to_sfixed(0.79,5,4),	to_sfixed(2.57,5,4),	to_sfixed(580,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.86,5,4),	to_sfixed(1.35,5,4),	to_sfixed(2.32,5,4),	to_sfixed(18,5,4),	to_sfixed(122,5,4),	to_sfixed(1.51,5,4),	to_sfixed(1.25,5,4),	to_sfixed(0.21,5,4),	to_sfixed(0.94,5,4),	to_sfixed(4.1,5,4),	to_sfixed(0.76,5,4),	to_sfixed(1.29,5,4),	to_sfixed(630,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.88,5,4),	to_sfixed(2.99,5,4),	to_sfixed(2.4,5,4),	to_sfixed(20,5,4),	to_sfixed(104,5,4),	to_sfixed(1.3,5,4),	to_sfixed(1.22,5,4),	to_sfixed(0.24,5,4),	to_sfixed(0.83,5,4),	to_sfixed(5.4,5,4),	to_sfixed(0.74,5,4),	to_sfixed(1.42,5,4),	to_sfixed(530,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.81,5,4),	to_sfixed(2.31,5,4),	to_sfixed(2.4,5,4),	to_sfixed(24,5,4),	to_sfixed(98,5,4),	to_sfixed(1.15,5,4),	to_sfixed(1.09,5,4),	to_sfixed(0.27,5,4),	to_sfixed(0.83,5,4),	to_sfixed(5.7,5,4),	to_sfixed(0.66,5,4),	to_sfixed(1.36,5,4),	to_sfixed(560,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.7,5,4),		to_sfixed(3.55,5,4),	to_sfixed(2.36,5,4),	to_sfixed(21.5,5,4),	to_sfixed(106,5,4),	to_sfixed(1.7,5,4),	to_sfixed(1.2,5,4),	to_sfixed(0.17,5,4),	to_sfixed(0.84,5,4),	to_sfixed(5,5,4),		to_sfixed(0.78,5,4),	to_sfixed(1.29,5,4),	to_sfixed(600,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.51,5,4),	to_sfixed(1.24,5,4),	to_sfixed(2.25,5,4),	to_sfixed(17.5,5,4),	to_sfixed(85,5,4),	to_sfixed(2,5,4),		to_sfixed(0.58,5,4),	to_sfixed(0.6,5,4),	to_sfixed(1.25,5,4),	to_sfixed(5.45,5,4),	to_sfixed(0.75,5,4),	to_sfixed(1.51,5,4),	to_sfixed(650,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.6,5,4),		to_sfixed(2.46,5,4),	to_sfixed(2.2,5,4),	to_sfixed(18.5,5,4),	to_sfixed(94,5,4),	to_sfixed(1.62,5,4),	to_sfixed(0.66,5,4),	to_sfixed(0.63,5,4),	to_sfixed(0.94,5,4),	to_sfixed(7.1,5,4),	to_sfixed(0.73,5,4),	to_sfixed(1.58,5,4),	to_sfixed(695,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.25,5,4),	to_sfixed(4.72,5,4),	to_sfixed(2.54,5,4),	to_sfixed(21,5,4),	to_sfixed(89,5,4),	to_sfixed(1.38,5,4),	to_sfixed(0.47,5,4),	to_sfixed(0.53,5,4),	to_sfixed(0.8,5,4),	to_sfixed(3.85,5,4),	to_sfixed(0.75,5,4),	to_sfixed(1.27,5,4),	to_sfixed(720,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.53,5,4),	to_sfixed(5.51,5,4),	to_sfixed(2.64,5,4),	to_sfixed(25,5,4),	to_sfixed(96,5,4),	to_sfixed(1.79,5,4),	to_sfixed(0.6,5,4),	to_sfixed(0.63,5,4),	to_sfixed(1.1,5,4),	to_sfixed(5,5,4),		to_sfixed(0.82,5,4),	to_sfixed(1.69,5,4),	to_sfixed(515,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.49,5,4),	to_sfixed(3.59,5,4),	to_sfixed(2.19,5,4),	to_sfixed(19.5,5,4),	to_sfixed(88,5,4),	to_sfixed(1.62,5,4),	to_sfixed(0.48,5,4),	to_sfixed(0.58,5,4),	to_sfixed(0.88,5,4),	to_sfixed(5.7,5,4),	to_sfixed(0.81,5,4),	to_sfixed(1.82,5,4),	to_sfixed(580,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.84,5,4),	to_sfixed(2.96,5,4),	to_sfixed(2.61,5,4),	to_sfixed(24,5,4),	to_sfixed(101,5,4),	to_sfixed(2.32,5,4),	to_sfixed(0.6,5,4),	to_sfixed(0.53,5,4),	to_sfixed(0.81,5,4),	to_sfixed(4.92,5,4),	to_sfixed(0.89,5,4),	to_sfixed(2.15,5,4),	to_sfixed(590,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.93,5,4),	to_sfixed(2.81,5,4),	to_sfixed(2.7,5,4),	to_sfixed(21,5,4),	to_sfixed(96,5,4),	to_sfixed(1.54,5,4),	to_sfixed(0.5,5,4),	to_sfixed(0.53,5,4),	to_sfixed(0.75,5,4),	to_sfixed(4.6,5,4),	to_sfixed(0.77,5,4),	to_sfixed(2.31,5,4),	to_sfixed(600,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.36,5,4),	to_sfixed(2.56,5,4),	to_sfixed(2.35,5,4),	to_sfixed(20,5,4),	to_sfixed(89,5,4),	to_sfixed(1.4,5,4),	to_sfixed(0.5,5,4),	to_sfixed(0.37,5,4),	to_sfixed(0.64,5,4),	to_sfixed(5.6,5,4),	to_sfixed(0.7,5,4),	to_sfixed(2.47,5,4),	to_sfixed(780,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.52,5,4),	to_sfixed(3.17,5,4),	to_sfixed(2.72,5,4),	to_sfixed(23.5,5,4),	to_sfixed(97,5,4),	to_sfixed(1.55,5,4),	to_sfixed(0.52,5,4),	to_sfixed(0.5,5,4),	to_sfixed(0.55,5,4),	to_sfixed(4.35,5,4),	to_sfixed(0.89,5,4),	to_sfixed(2.06,5,4),	to_sfixed(520,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.62,5,4),	to_sfixed(4.95,5,4),	to_sfixed(2.35,5,4),	to_sfixed(20,5,4),	to_sfixed(92,5,4),	to_sfixed(2,5,4),		to_sfixed(0.8,5,4),	to_sfixed(0.47,5,4),	to_sfixed(1.02,5,4),	to_sfixed(4.4,5,4),	to_sfixed(0.91,5,4),	to_sfixed(2.05,5,4),	to_sfixed(550,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.25,5,4),	to_sfixed(3.88,5,4),	to_sfixed(2.2,5,4),	to_sfixed(18.5,5,4),	to_sfixed(112,5,4),	to_sfixed(1.38,5,4),	to_sfixed(0.78,5,4),	to_sfixed(0.29,5,4),	to_sfixed(1.14,5,4),	to_sfixed(8.21,5,4),	to_sfixed(0.65,5,4),	to_sfixed(2,5,4),		to_sfixed(855,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.16,5,4),	to_sfixed(3.57,5,4),	to_sfixed(2.15,5,4),	to_sfixed(21,5,4),	to_sfixed(102,5,4),	to_sfixed(1.5,5,4),	to_sfixed(0.55,5,4),	to_sfixed(0.43,5,4),	to_sfixed(1.3,5,4),	to_sfixed(4,5,4),		to_sfixed(0.6,5,4),	to_sfixed(1.68,5,4),	to_sfixed(830,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.88,5,4),	to_sfixed(5.04,5,4),	to_sfixed(2.23,5,4),	to_sfixed(20,5,4),	to_sfixed(80,5,4),	to_sfixed(0.98,5,4),	to_sfixed(0.34,5,4),	to_sfixed(0.4,5,4),	to_sfixed(0.68,5,4),	to_sfixed(4.9,5,4),	to_sfixed(0.58,5,4),	to_sfixed(1.33,5,4),	to_sfixed(415,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.87,5,4),	to_sfixed(4.61,5,4),	to_sfixed(2.48,5,4),	to_sfixed(21.5,5,4),	to_sfixed(86,5,4),	to_sfixed(1.7,5,4),	to_sfixed(0.65,5,4),	to_sfixed(0.47,5,4),	to_sfixed(0.86,5,4),	to_sfixed(7.65,5,4),	to_sfixed(0.54,5,4),	to_sfixed(1.86,5,4),	to_sfixed(625,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.32,5,4),	to_sfixed(3.24,5,4),	to_sfixed(2.38,5,4),	to_sfixed(21.5,5,4),	to_sfixed(92,5,4),	to_sfixed(1.93,5,4),	to_sfixed(0.76,5,4),	to_sfixed(0.45,5,4),	to_sfixed(1.25,5,4),	to_sfixed(8.42,5,4),	to_sfixed(0.55,5,4),	to_sfixed(1.62,5,4),	to_sfixed(650,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.08,5,4),	to_sfixed(3.9,5,4),	to_sfixed(2.36,5,4),	to_sfixed(21.5,5,4),	to_sfixed(113,5,4),	to_sfixed(1.41,5,4),	to_sfixed(1.39,5,4),	to_sfixed(0.34,5,4),	to_sfixed(1.14,5,4),	to_sfixed(9.40,5,4),	to_sfixed(0.57,5,4),	to_sfixed(1.33,5,4),	to_sfixed(550,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.5,5,4),		to_sfixed(3.12,5,4),	to_sfixed(2.62,5,4),	to_sfixed(24,5,4),	to_sfixed(123,5,4),	to_sfixed(1.4,5,4),	to_sfixed(1.57,5,4),	to_sfixed(0.22,5,4),	to_sfixed(1.25,5,4),	to_sfixed(8.60,5,4),	to_sfixed(0.59,5,4),	to_sfixed(1.3,5,4),	to_sfixed(500,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.79,5,4),	to_sfixed(2.67,5,4),	to_sfixed(2.48,5,4),	to_sfixed(22,5,4),	to_sfixed(112,5,4),	to_sfixed(1.48,5,4),	to_sfixed(1.36,5,4),	to_sfixed(0.24,5,4),	to_sfixed(1.26,5,4),	to_sfixed(10.8,5,4),	to_sfixed(0.48,5,4),	to_sfixed(1.47,5,4),	to_sfixed(480,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.11,5,4),	to_sfixed(1.9,5,4),	to_sfixed(2.75,5,4),	to_sfixed(25.5,5,4),	to_sfixed(116,5,4),	to_sfixed(2.2,5,4),	to_sfixed(1.28,5,4),	to_sfixed(0.26,5,4),	to_sfixed(1.56,5,4),	to_sfixed(7.1,5,4),	to_sfixed(0.61,5,4),	to_sfixed(1.33,5,4),	to_sfixed(425,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.23,5,4),	to_sfixed(3.3,5,4),	to_sfixed(2.28,5,4),	to_sfixed(18.5,5,4),	to_sfixed(98,5,4),	to_sfixed(1.8,5,4),	to_sfixed(0.83,5,4),	to_sfixed(0.61,5,4),	to_sfixed(1.87,5,4),	to_sfixed(10.52,5,4),to_sfixed(0.56,5,4),	to_sfixed(1.51,5,4),	to_sfixed(675,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.58,5,4),	to_sfixed(1.29,5,4),	to_sfixed(2.1,5,4),	to_sfixed(20,5,4),	to_sfixed(103,5,4),	to_sfixed(1.48,5,4),	to_sfixed(0.58,5,4),	to_sfixed(0.53,5,4),	to_sfixed(1.4,5,4),	to_sfixed(7.6,5,4),	to_sfixed(0.58,5,4),	to_sfixed(1.55,5,4),	to_sfixed(640,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.17,5,4),	to_sfixed(5.19,5,4),	to_sfixed(2.32,5,4),	to_sfixed(22,5,4),	to_sfixed(93,5,4),	to_sfixed(1.74,5,4),	to_sfixed(0.63,5,4),	to_sfixed(0.61,5,4),	to_sfixed(1.55,5,4),	to_sfixed(7.9,5,4),	to_sfixed(0.6,5,4),	to_sfixed(1.48,5,4),	to_sfixed(725,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.84,5,4),	to_sfixed(4.12,5,4),	to_sfixed(2.38,5,4),	to_sfixed(19.5,5,4),	to_sfixed(89,5,4),	to_sfixed(1.8,5,4),	to_sfixed(0.83,5,4),	to_sfixed(0.48,5,4),	to_sfixed(1.56,5,4),	to_sfixed(9.01,5,4),	to_sfixed(0.57,5,4),	to_sfixed(1.64,5,4),	to_sfixed(480,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.45,5,4),	to_sfixed(3.03,5,4),	to_sfixed(2.64,5,4),	to_sfixed(27,5,4),	to_sfixed(97,5,4),	to_sfixed(1.9,5,4),	to_sfixed(0.58,5,4),	to_sfixed(0.63,5,4),	to_sfixed(1.14,5,4),	to_sfixed(7.5,5,4),	to_sfixed(0.67,5,4),	to_sfixed(1.73,5,4),	to_sfixed(880,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(14.34,5,4),	to_sfixed(1.68,5,4),	to_sfixed(2.7,5,4),	to_sfixed(25,5,4),	to_sfixed(98,5,4),	to_sfixed(2.8,5,4),	to_sfixed(1.31,5,4),	to_sfixed(0.53,5,4),	to_sfixed(2.7,5,4),	to_sfixed(13,5,4),	to_sfixed(0.57,5,4),	to_sfixed(1.96,5,4),	to_sfixed(660,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.48,5,4),	to_sfixed(1.67,5,4),	to_sfixed(2.64,5,4),	to_sfixed(22.5,5,4),	to_sfixed(89,5,4),	to_sfixed(2.6,5,4),	to_sfixed(1.1,5,4),	to_sfixed(0.52,5,4),	to_sfixed(2.29,5,4),	to_sfixed(11.75,5,4),to_sfixed(0.57,5,4),	to_sfixed(1.78,5,4),	to_sfixed(620,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.36,5,4),	to_sfixed(3.83,5,4),	to_sfixed(2.38,5,4),	to_sfixed(21,5,4),	to_sfixed(88,5,4),	to_sfixed(2.3,5,4),	to_sfixed(0.92,5,4),	to_sfixed(0.5,5,4),	to_sfixed(1.04,5,4),	to_sfixed(7.65,5,4),	to_sfixed(0.56,5,4),	to_sfixed(1.58,5,4),	to_sfixed(520,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.69,5,4),	to_sfixed(3.26,5,4),	to_sfixed(2.54,5,4),	to_sfixed(20,5,4),	to_sfixed(107,5,4),	to_sfixed(1.83,5,4),	to_sfixed(0.56,5,4),	to_sfixed(0.5,5,4),	to_sfixed(0.8,5,4),	to_sfixed(5.88,5,4),	to_sfixed(0.96,5,4),	to_sfixed(1.82,5,4),	to_sfixed(680,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.85,5,4),	to_sfixed(3.27,5,4),	to_sfixed(2.58,5,4),	to_sfixed(22,5,4),	to_sfixed(106,5,4),	to_sfixed(1.65,5,4),	to_sfixed(0.6,5,4),	to_sfixed(0.6,5,4),	to_sfixed(0.96,5,4),	to_sfixed(5.58,5,4),	to_sfixed(0.87,5,4),	to_sfixed(2.11,5,4),	to_sfixed(570,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.96,5,4),	to_sfixed(3.45,5,4),	to_sfixed(2.35,5,4),	to_sfixed(18.5,5,4),	to_sfixed(106,5,4),	to_sfixed(1.39,5,4),	to_sfixed(0.7,5,4),	to_sfixed(0.4,5,4),	to_sfixed(0.94,5,4),	to_sfixed(5.28,5,4),	to_sfixed(0.68,5,4),	to_sfixed(1.75,5,4),	to_sfixed(675,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.78,5,4),	to_sfixed(2.76,5,4),	to_sfixed(2.3,5,4),	to_sfixed(22,5,4),	to_sfixed(90,5,4),	to_sfixed(1.35,5,4),	to_sfixed(0.68,5,4),	to_sfixed(0.41,5,4),	to_sfixed(1.03,5,4),	to_sfixed(9.58,5,4),	to_sfixed(0.7,5,4),	to_sfixed(1.68,5,4),	to_sfixed(615,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.73,5,4),	to_sfixed(4.36,5,4),	to_sfixed(2.26,5,4),	to_sfixed(22.5,5,4),	to_sfixed(88,5,4),	to_sfixed(1.28,5,4),	to_sfixed(0.47,5,4),	to_sfixed(0.52,5,4),	to_sfixed(1.15,5,4),	to_sfixed(6.62,5,4),	to_sfixed(0.78,5,4),	to_sfixed(1.75,5,4),	to_sfixed(520,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.45,5,4),	to_sfixed(3.7,5,4),	to_sfixed(2.6,5,4),	to_sfixed(23,5,4),	to_sfixed(111,5,4),	to_sfixed(1.7,5,4),	to_sfixed(0.92,5,4),	to_sfixed(0.43,5,4),	to_sfixed(1.46,5,4),	to_sfixed(10.68,5,4),to_sfixed(0.85,5,4),	to_sfixed(1.56,5,4),	to_sfixed(695,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.82,5,4),	to_sfixed(3.37,5,4),	to_sfixed(2.3,5,4),	to_sfixed(19.5,5,4),	to_sfixed(88,5,4),	to_sfixed(1.48,5,4),	to_sfixed(0.66,5,4),	to_sfixed(0.4,5,4),	to_sfixed(0.97,5,4),	to_sfixed(10.26,5,4),to_sfixed(0.72,5,4),	to_sfixed(1.75,5,4),	to_sfixed(685,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.58,5,4),	to_sfixed(2.58,5,4),	to_sfixed(2.69,5,4),	to_sfixed(24.5,5,4),	to_sfixed(105,5,4),	to_sfixed(1.55,5,4),	to_sfixed(0.84,5,4),	to_sfixed(0.39,5,4),	to_sfixed(1.54,5,4),	to_sfixed(8.66,5,4),	to_sfixed(0.74,5,4),	to_sfixed(1.8,5,4),	to_sfixed(750,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.4,5,4),		to_sfixed(4.6,5,4),	to_sfixed(2.86,5,4),	to_sfixed(25,5,4),	to_sfixed(112,5,4),	to_sfixed(1.98,5,4),	to_sfixed(0.96,5,4),	to_sfixed(0.27,5,4),	to_sfixed(1.11,5,4),	to_sfixed(8.5,5,4),	to_sfixed(0.67,5,4),	to_sfixed(1.92,5,4),	to_sfixed(630,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.2,5,4),		to_sfixed(3.03,5,4),	to_sfixed(2.32,5,4),	to_sfixed(19,5,4),	to_sfixed(96,5,4),	to_sfixed(1.25,5,4),	to_sfixed(0.49,5,4),	to_sfixed(0.4,5,4),	to_sfixed(0.73,5,4),	to_sfixed(5.5,5,4),	to_sfixed(0.66,5,4),	to_sfixed(1.83,5,4),	to_sfixed(510,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(12.77,5,4),	to_sfixed(2.39,5,4),	to_sfixed(2.28,5,4),	to_sfixed(19.5,5,4),	to_sfixed(86,5,4),	to_sfixed(1.39,5,4),	to_sfixed(0.51,5,4),	to_sfixed(0.48,5,4),	to_sfixed(0.64,5,4),	to_sfixed(9.90,5,4),	to_sfixed(0.57,5,4),	to_sfixed(1.63,5,4),	to_sfixed(470,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(14.16,5,4),	to_sfixed(2.51,5,4),	to_sfixed(2.48,5,4),	to_sfixed(20,5,4),	to_sfixed(91,5,4),	to_sfixed(1.68,5,4),	to_sfixed(0.7,5,4),	to_sfixed(0.44,5,4),	to_sfixed(1.24,5,4),	to_sfixed(9.7,5,4),	to_sfixed(0.62,5,4),	to_sfixed(1.71,5,4),	to_sfixed(660,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.71,5,4),	to_sfixed(5.65,5,4),	to_sfixed(2.45,5,4),	to_sfixed(20.5,5,4),	to_sfixed(95,5,4),	to_sfixed(1.68,5,4),	to_sfixed(0.61,5,4),	to_sfixed(0.52,5,4),	to_sfixed(1.06,5,4),	to_sfixed(7.7,5,4),	to_sfixed(0.64,5,4),	to_sfixed(1.74,5,4),	to_sfixed(740,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.4,5,4),		to_sfixed(3.91,5,4),	to_sfixed(2.48,5,4),	to_sfixed(23,5,4),	to_sfixed(102,5,4),	to_sfixed(1.8,5,4),	to_sfixed(0.75,5,4),	to_sfixed(0.43,5,4),	to_sfixed(1.41,5,4),	to_sfixed(7.3,5,4),	to_sfixed(0.7,5,4),	to_sfixed(1.56,5,4),	to_sfixed(750,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.27,5,4),	to_sfixed(4.28,5,4),	to_sfixed(2.26,5,4),	to_sfixed(20,5,4),	to_sfixed(120,5,4),	to_sfixed(1.59,5,4),	to_sfixed(0.69,5,4),	to_sfixed(0.43,5,4),	to_sfixed(1.35,5,4),	to_sfixed(10.2,5,4),	to_sfixed(0.59,5,4),	to_sfixed(1.56,5,4),	to_sfixed(835,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(13.17,5,4),	to_sfixed(2.59,5,4),	to_sfixed(2.37,5,4),	to_sfixed(20,5,4),	to_sfixed(120,5,4),	to_sfixed(1.65,5,4),	to_sfixed(0.68,5,4),	to_sfixed(0.53,5,4),	to_sfixed(1.46,5,4),	to_sfixed(9.3,5,4),	to_sfixed(0.6,5,4),	to_sfixed(1.62,5,4),	to_sfixed(840,5,4)),
		(to_sfixed(3,5,4),	to_sfixed(14.13,5,4),	to_sfixed(4.1,5,4),	to_sfixed(2.74,5,4),	to_sfixed(24.5,5,4),	to_sfixed(96,5,4),	to_sfixed(2.05,5,4),	to_sfixed(0.76,5,4),	to_sfixed(0.56,5,4),	to_sfixed(1.35,5,4),	to_sfixed(9.2,5,4),	to_sfixed(0.61,5,4),	to_sfixed(1.6,5,4),	to_sfixed(560,5,4))
	); 
	
end package body;

    