--=============================================================================
--    This file is part of FPGA_NEURAL-Network.
--
--    FPGA_NEURAL-Network is free software: you can redistribute it and/or 
--    modify it under the terms of the GNU General Public License as published 
--    by the Free Software Foundation, either version 3 of the License, or
--    (at your option) any later version.
--
--    FPGA_NEURAL-Network is distributed in the hope that it will be useful,
--    but WITHOUT ANY WARRANTY; without even the implied warranty of
--    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--    GNU General Public License for more details.
--
--    You should have received a copy of the GNU General Public License
--    along with FPGA_NEURAL-Network.  
--		if not, see <http://www.gnu.org/licenses/>.

--=============================================================================
--	FILE NAME			: INPUT_ROM.vhd
--	PROJECT				: FPGA_NEURAL-Network
--	ENTITY				: INPUT_ROM
--	ARCHITECTURE		: rtl
--=============================================================================
--	AUTORS(s)			: Agostini, N;
--	DEPARTMENT      	: Electrical Engineering (UFRGS)
--	DATE					: Dec 14, 2014
--=============================================================================
--	Description:
--	
--=============================================================================

library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all; -- is the to unsigned really required????
	use work.fixed_pkg.all; -- ieee_proposed for compatibility version
	use work.NN_TYPES_pkg.all;
	use work.INPUT_ROM_pkg.all;

--=============================================================================
-- Entity declaration for INPUT_ROM
--=============================================================================
entity INPUT_ROM is 
	port (
		clk				:	in std_logic;
		SAMPLE_NUMBER 	: 	in std_logic_vector (7 downto 0);
		SELECTED_INPUT	: 	out ARRAY_OF_SFIXED
	);
end INPUT_ROM;

--=============================================================================
-- architecture declaration
--=============================================================================
architecture RTL of INPUT_ROM is
-- Constants
	constant INPUTS_TABLE : INPUT_TABLE(0 to SAMPLE_SIZE-1) := (
					(to_sfixed(0.9595,1,L_SIZE), to_sfixed(0.2948,1,L_SIZE), to_sfixed(0.7523,1,L_SIZE), to_sfixed(0.5200,1,L_SIZE), to_sfixed(0.7840,1,L_SIZE), to_sfixed(0.7216,1,L_SIZE), to_sfixed(0.6024,1,L_SIZE), to_sfixed(0.4242,1,L_SIZE), to_sfixed(0.6397,1,L_SIZE), to_sfixed(0.4338,1,L_SIZE), to_sfixed(0.6082,1,L_SIZE), to_sfixed(0.9800,1,L_SIZE), to_sfixed(0.6339,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8901,1,L_SIZE), to_sfixed(0.3069,1,L_SIZE), to_sfixed(0.6625,1,L_SIZE), to_sfixed(0.3733,1,L_SIZE), to_sfixed(0.6173,1,L_SIZE), to_sfixed(0.6830,1,L_SIZE), to_sfixed(0.5433,1,L_SIZE), to_sfixed(0.3939,1,L_SIZE), to_sfixed(0.3575,1,L_SIZE), to_sfixed(0.3369,1,L_SIZE), to_sfixed(0.6140,1,L_SIZE), to_sfixed(0.8500,1,L_SIZE), to_sfixed(0.6250,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8874,1,L_SIZE), to_sfixed(0.4069,1,L_SIZE), to_sfixed(0.8266,1,L_SIZE), to_sfixed(0.6200,1,L_SIZE), to_sfixed(0.6235,1,L_SIZE), to_sfixed(0.7216,1,L_SIZE), to_sfixed(0.6378,1,L_SIZE), to_sfixed(0.4545,1,L_SIZE), to_sfixed(0.7849,1,L_SIZE), to_sfixed(0.4369,1,L_SIZE), to_sfixed(0.6023,1,L_SIZE), to_sfixed(0.7925,1,L_SIZE), to_sfixed(0.7054,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9690,1,L_SIZE), to_sfixed(0.3362,1,L_SIZE), to_sfixed(0.7740,1,L_SIZE), to_sfixed(0.5600,1,L_SIZE), to_sfixed(0.6975,1,L_SIZE), to_sfixed(0.9923,1,L_SIZE), to_sfixed(0.6870,1,L_SIZE), to_sfixed(0.3636,1,L_SIZE), to_sfixed(0.6089,1,L_SIZE), to_sfixed(0.6000,1,L_SIZE), to_sfixed(0.5029,1,L_SIZE), to_sfixed(0.8625,1,L_SIZE), to_sfixed(0.8810,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8928,1,L_SIZE), to_sfixed(0.4466,1,L_SIZE), to_sfixed(0.8885,1,L_SIZE), to_sfixed(0.7000,1,L_SIZE), to_sfixed(0.7284,1,L_SIZE), to_sfixed(0.7216,1,L_SIZE), to_sfixed(0.5295,1,L_SIZE), to_sfixed(0.5909,1,L_SIZE), to_sfixed(0.5084,1,L_SIZE), to_sfixed(0.3323,1,L_SIZE), to_sfixed(0.6082,1,L_SIZE), to_sfixed(0.7325,1,L_SIZE), to_sfixed(0.4375,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9575,1,L_SIZE), to_sfixed(0.3034,1,L_SIZE), to_sfixed(0.7585,1,L_SIZE), to_sfixed(0.5067,1,L_SIZE), to_sfixed(0.6914,1,L_SIZE), to_sfixed(0.8428,1,L_SIZE), to_sfixed(0.6673,1,L_SIZE), to_sfixed(0.5152,1,L_SIZE), to_sfixed(0.5503,1,L_SIZE), to_sfixed(0.5192,1,L_SIZE), to_sfixed(0.6140,1,L_SIZE), to_sfixed(0.7125,1,L_SIZE), to_sfixed(0.8631,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9703,1,L_SIZE), to_sfixed(0.3224,1,L_SIZE), to_sfixed(0.7585,1,L_SIZE), to_sfixed(0.4867,1,L_SIZE), to_sfixed(0.5926,1,L_SIZE), to_sfixed(0.6443,1,L_SIZE), to_sfixed(0.4961,1,L_SIZE), to_sfixed(0.4545,1,L_SIZE), to_sfixed(0.5531,1,L_SIZE), to_sfixed(0.4038,1,L_SIZE), to_sfixed(0.5965,1,L_SIZE), to_sfixed(0.8950,1,L_SIZE), to_sfixed(0.7679,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9481,1,L_SIZE), to_sfixed(0.3707,1,L_SIZE), to_sfixed(0.8080,1,L_SIZE), to_sfixed(0.5867,1,L_SIZE), to_sfixed(0.7469,1,L_SIZE), to_sfixed(0.6701,1,L_SIZE), to_sfixed(0.4941,1,L_SIZE), to_sfixed(0.4697,1,L_SIZE), to_sfixed(0.3492,1,L_SIZE), to_sfixed(0.3885,1,L_SIZE), to_sfixed(0.6199,1,L_SIZE), to_sfixed(0.8950,1,L_SIZE), to_sfixed(0.7708,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.2828,1,L_SIZE), to_sfixed(0.6718,1,L_SIZE), to_sfixed(0.4667,1,L_SIZE), to_sfixed(0.5988,1,L_SIZE), to_sfixed(0.7216,1,L_SIZE), to_sfixed(0.5866,1,L_SIZE), to_sfixed(0.4394,1,L_SIZE), to_sfixed(0.5531,1,L_SIZE), to_sfixed(0.4000,1,L_SIZE), to_sfixed(0.6316,1,L_SIZE), to_sfixed(0.7125,1,L_SIZE), to_sfixed(0.6220,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9346,1,L_SIZE), to_sfixed(0.2328,1,L_SIZE), to_sfixed(0.7028,1,L_SIZE), to_sfixed(0.5333,1,L_SIZE), to_sfixed(0.6049,1,L_SIZE), to_sfixed(0.7680,1,L_SIZE), to_sfixed(0.6201,1,L_SIZE), to_sfixed(0.3333,1,L_SIZE), to_sfixed(0.5168,1,L_SIZE), to_sfixed(0.5554,1,L_SIZE), to_sfixed(0.5906,1,L_SIZE), to_sfixed(0.8875,1,L_SIZE), to_sfixed(0.6220,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9508,1,L_SIZE), to_sfixed(0.3724,1,L_SIZE), to_sfixed(0.7121,1,L_SIZE), to_sfixed(0.6000,1,L_SIZE), to_sfixed(0.6481,1,L_SIZE), to_sfixed(0.7603,1,L_SIZE), to_sfixed(0.6535,1,L_SIZE), to_sfixed(0.3333,1,L_SIZE), to_sfixed(0.6648,1,L_SIZE), to_sfixed(0.4423,1,L_SIZE), to_sfixed(0.7310,1,L_SIZE), to_sfixed(0.7925,1,L_SIZE), to_sfixed(0.8988,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9521,1,L_SIZE), to_sfixed(0.2552,1,L_SIZE), to_sfixed(0.7183,1,L_SIZE), to_sfixed(0.5600,1,L_SIZE), to_sfixed(0.5864,1,L_SIZE), to_sfixed(0.5670,1,L_SIZE), to_sfixed(0.4783,1,L_SIZE), to_sfixed(0.3939,1,L_SIZE), to_sfixed(0.4385,1,L_SIZE), to_sfixed(0.3846,1,L_SIZE), to_sfixed(0.6842,1,L_SIZE), to_sfixed(0.7050,1,L_SIZE), to_sfixed(0.7619,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9272,1,L_SIZE), to_sfixed(0.2983,1,L_SIZE), to_sfixed(0.7461,1,L_SIZE), to_sfixed(0.5333,1,L_SIZE), to_sfixed(0.5494,1,L_SIZE), to_sfixed(0.6701,1,L_SIZE), to_sfixed(0.5433,1,L_SIZE), to_sfixed(0.4394,1,L_SIZE), to_sfixed(0.5056,1,L_SIZE), to_sfixed(0.4308,1,L_SIZE), to_sfixed(0.6725,1,L_SIZE), to_sfixed(0.7250,1,L_SIZE), to_sfixed(0.7857,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9946,1,L_SIZE), to_sfixed(0.2983,1,L_SIZE), to_sfixed(0.7399,1,L_SIZE), to_sfixed(0.3800,1,L_SIZE), to_sfixed(0.5617,1,L_SIZE), to_sfixed(0.7990,1,L_SIZE), to_sfixed(0.7264,1,L_SIZE), to_sfixed(0.6515,1,L_SIZE), to_sfixed(0.7849,1,L_SIZE), to_sfixed(0.4154,1,L_SIZE), to_sfixed(0.7310,1,L_SIZE), to_sfixed(0.6825,1,L_SIZE), to_sfixed(0.6845,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9697,1,L_SIZE), to_sfixed(0.3224,1,L_SIZE), to_sfixed(0.7368,1,L_SIZE), to_sfixed(0.4000,1,L_SIZE), to_sfixed(0.6296,1,L_SIZE), to_sfixed(0.8505,1,L_SIZE), to_sfixed(0.7165,1,L_SIZE), to_sfixed(0.4394,1,L_SIZE), to_sfixed(0.8268,1,L_SIZE), to_sfixed(0.5769,1,L_SIZE), to_sfixed(0.7018,1,L_SIZE), to_sfixed(0.7500,1,L_SIZE), to_sfixed(0.9208,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9191,1,L_SIZE), to_sfixed(0.3121,1,L_SIZE), to_sfixed(0.8359,1,L_SIZE), to_sfixed(0.5733,1,L_SIZE), to_sfixed(0.6914,1,L_SIZE), to_sfixed(0.7345,1,L_SIZE), to_sfixed(0.5728,1,L_SIZE), to_sfixed(0.4545,1,L_SIZE), to_sfixed(0.4078,1,L_SIZE), to_sfixed(0.5615,1,L_SIZE), to_sfixed(0.7485,1,L_SIZE), to_sfixed(0.7200,1,L_SIZE), to_sfixed(0.7798,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9643,1,L_SIZE), to_sfixed(0.3310,1,L_SIZE), to_sfixed(0.8421,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(0.7407,1,L_SIZE), to_sfixed(0.7216,1,L_SIZE), to_sfixed(0.6181,1,L_SIZE), to_sfixed(0.5000,1,L_SIZE), to_sfixed(0.5503,1,L_SIZE), to_sfixed(0.4769,1,L_SIZE), to_sfixed(0.6257,1,L_SIZE), to_sfixed(0.6625,1,L_SIZE), to_sfixed(0.7619,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9326,1,L_SIZE), to_sfixed(0.2707,1,L_SIZE), to_sfixed(0.8111,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(0.7099,1,L_SIZE), to_sfixed(0.7603,1,L_SIZE), to_sfixed(0.6693,1,L_SIZE), to_sfixed(0.6061,1,L_SIZE), to_sfixed(0.4804,1,L_SIZE), to_sfixed(0.5077,1,L_SIZE), to_sfixed(0.6608,1,L_SIZE), to_sfixed(0.6425,1,L_SIZE), to_sfixed(0.6726,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9568,1,L_SIZE), to_sfixed(0.2741,1,L_SIZE), to_sfixed(0.7678,1,L_SIZE), to_sfixed(0.5500,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(0.8505,1,L_SIZE), to_sfixed(0.7736,1,L_SIZE), to_sfixed(0.4848,1,L_SIZE), to_sfixed(0.5196,1,L_SIZE), to_sfixed(0.6692,1,L_SIZE), to_sfixed(0.7193,1,L_SIZE), to_sfixed(0.7050,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9198,1,L_SIZE), to_sfixed(0.5345,1,L_SIZE), to_sfixed(0.7926,1,L_SIZE), to_sfixed(0.5067,1,L_SIZE), to_sfixed(0.7160,1,L_SIZE), to_sfixed(0.6959,1,L_SIZE), to_sfixed(0.5965,1,L_SIZE), to_sfixed(0.2576,1,L_SIZE), to_sfixed(0.4637,1,L_SIZE), to_sfixed(0.3923,1,L_SIZE), to_sfixed(0.5614,1,L_SIZE), to_sfixed(0.8400,1,L_SIZE), to_sfixed(0.5030,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9481,1,L_SIZE), to_sfixed(0.2810,1,L_SIZE), to_sfixed(0.7059,1,L_SIZE), to_sfixed(0.5333,1,L_SIZE), to_sfixed(0.7778,1,L_SIZE), to_sfixed(0.7732,1,L_SIZE), to_sfixed(0.6240,1,L_SIZE), to_sfixed(0.3636,1,L_SIZE), to_sfixed(0.5866,1,L_SIZE), to_sfixed(0.4346,1,L_SIZE), to_sfixed(0.6374,1,L_SIZE), to_sfixed(0.9275,1,L_SIZE), to_sfixed(0.4643,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8719,1,L_SIZE), to_sfixed(0.6552,1,L_SIZE), to_sfixed(0.8204,1,L_SIZE), to_sfixed(0.6200,1,L_SIZE), to_sfixed(0.6296,1,L_SIZE), to_sfixed(0.6211,1,L_SIZE), to_sfixed(0.4744,1,L_SIZE), to_sfixed(0.3788,1,L_SIZE), to_sfixed(0.5531,1,L_SIZE), to_sfixed(0.3462,1,L_SIZE), to_sfixed(0.6023,1,L_SIZE), to_sfixed(0.8800,1,L_SIZE), to_sfixed(0.4583,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9245,1,L_SIZE), to_sfixed(0.3207,1,L_SIZE), to_sfixed(0.7307,1,L_SIZE), to_sfixed(0.5533,1,L_SIZE), to_sfixed(0.6235,1,L_SIZE), to_sfixed(0.6727,1,L_SIZE), to_sfixed(0.5669,1,L_SIZE), to_sfixed(0.4091,1,L_SIZE), to_sfixed(0.4721,1,L_SIZE), to_sfixed(0.2923,1,L_SIZE), to_sfixed(0.6491,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.6161,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8665,1,L_SIZE), to_sfixed(0.2759,1,L_SIZE), to_sfixed(0.7802,1,L_SIZE), to_sfixed(0.5933,1,L_SIZE), to_sfixed(0.5864,1,L_SIZE), to_sfixed(0.6392,1,L_SIZE), to_sfixed(0.4665,1,L_SIZE), to_sfixed(0.3939,1,L_SIZE), to_sfixed(0.4078,1,L_SIZE), to_sfixed(0.3023,1,L_SIZE), to_sfixed(0.6374,1,L_SIZE), to_sfixed(0.9075,1,L_SIZE), to_sfixed(0.6042,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9103,1,L_SIZE), to_sfixed(0.3121,1,L_SIZE), to_sfixed(0.8080,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(0.5926,1,L_SIZE), to_sfixed(0.6521,1,L_SIZE), to_sfixed(0.5138,1,L_SIZE), to_sfixed(0.4242,1,L_SIZE), to_sfixed(0.4637,1,L_SIZE), to_sfixed(0.2708,1,L_SIZE), to_sfixed(0.6550,1,L_SIZE), to_sfixed(0.9550,1,L_SIZE), to_sfixed(0.5030,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8800,1,L_SIZE), to_sfixed(0.3534,1,L_SIZE), to_sfixed(0.9969,1,L_SIZE), to_sfixed(0.8333,1,L_SIZE), to_sfixed(0.7654,1,L_SIZE), to_sfixed(0.6778,1,L_SIZE), to_sfixed(0.5276,1,L_SIZE), to_sfixed(0.7121,1,L_SIZE), to_sfixed(0.5363,1,L_SIZE), to_sfixed(0.2754,1,L_SIZE), to_sfixed(0.6608,1,L_SIZE), to_sfixed(0.8000,1,L_SIZE), to_sfixed(0.4940,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9029,1,L_SIZE), to_sfixed(0.3052,1,L_SIZE), to_sfixed(0.8111,1,L_SIZE), to_sfixed(0.5367,1,L_SIZE), to_sfixed(0.5741,1,L_SIZE), to_sfixed(0.7345,1,L_SIZE), to_sfixed(0.5787,1,L_SIZE), to_sfixed(0.5152,1,L_SIZE), to_sfixed(0.4050,1,L_SIZE), to_sfixed(0.3692,1,L_SIZE), to_sfixed(0.5380,1,L_SIZE), to_sfixed(0.8050,1,L_SIZE), to_sfixed(0.7113,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8968,1,L_SIZE), to_sfixed(0.2966,1,L_SIZE), to_sfixed(0.6625,1,L_SIZE), to_sfixed(0.5667,1,L_SIZE), to_sfixed(0.5802,1,L_SIZE), to_sfixed(0.6186,1,L_SIZE), to_sfixed(0.4311,1,L_SIZE), to_sfixed(0.4091,1,L_SIZE), to_sfixed(0.3771,1,L_SIZE), to_sfixed(0.3038,1,L_SIZE), to_sfixed(0.5965,1,L_SIZE), to_sfixed(0.6925,1,L_SIZE), to_sfixed(0.7649,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9353,1,L_SIZE), to_sfixed(0.3276,1,L_SIZE), to_sfixed(0.8669,1,L_SIZE), to_sfixed(0.6467,1,L_SIZE), to_sfixed(0.6605,1,L_SIZE), to_sfixed(0.7603,1,L_SIZE), to_sfixed(0.5846,1,L_SIZE), to_sfixed(0.5606,1,L_SIZE), to_sfixed(0.4916,1,L_SIZE), to_sfixed(0.3462,1,L_SIZE), to_sfixed(0.7310,1,L_SIZE), to_sfixed(0.8500,1,L_SIZE), to_sfixed(0.5446,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9454,1,L_SIZE), to_sfixed(0.2897,1,L_SIZE), to_sfixed(0.6842,1,L_SIZE), to_sfixed(0.5333,1,L_SIZE), to_sfixed(0.5926,1,L_SIZE), to_sfixed(0.6830,1,L_SIZE), to_sfixed(0.4587,1,L_SIZE), to_sfixed(0.3939,1,L_SIZE), to_sfixed(0.5531,1,L_SIZE), to_sfixed(0.3615,1,L_SIZE), to_sfixed(0.6082,1,L_SIZE), to_sfixed(0.8975,1,L_SIZE), to_sfixed(0.6161,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9258,1,L_SIZE), to_sfixed(0.2586,1,L_SIZE), to_sfixed(0.8359,1,L_SIZE), to_sfixed(0.7500,1,L_SIZE), to_sfixed(0.6235,1,L_SIZE), to_sfixed(0.7732,1,L_SIZE), to_sfixed(0.6398,1,L_SIZE), to_sfixed(0.4394,1,L_SIZE), to_sfixed(0.6648,1,L_SIZE), to_sfixed(0.4385,1,L_SIZE), to_sfixed(0.6959,1,L_SIZE), to_sfixed(0.6775,1,L_SIZE), to_sfixed(0.7649,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9157,1,L_SIZE), to_sfixed(0.2862,1,L_SIZE), to_sfixed(0.7307,1,L_SIZE), to_sfixed(0.6367,1,L_SIZE), to_sfixed(0.6543,1,L_SIZE), to_sfixed(0.7371,1,L_SIZE), to_sfixed(0.6280,1,L_SIZE), to_sfixed(0.3333,1,L_SIZE), to_sfixed(0.5447,1,L_SIZE), to_sfixed(0.5308,1,L_SIZE), to_sfixed(0.6374,1,L_SIZE), to_sfixed(0.7200,1,L_SIZE), to_sfixed(0.9018,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9225,1,L_SIZE), to_sfixed(0.3155,1,L_SIZE), to_sfixed(0.7307,1,L_SIZE), to_sfixed(0.5733,1,L_SIZE), to_sfixed(0.6420,1,L_SIZE), to_sfixed(0.6237,1,L_SIZE), to_sfixed(0.5295,1,L_SIZE), to_sfixed(0.6364,1,L_SIZE), to_sfixed(0.5503,1,L_SIZE), to_sfixed(0.2954,1,L_SIZE), to_sfixed(0.7193,1,L_SIZE), to_sfixed(0.7175,1,L_SIZE), to_sfixed(0.5893,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9278,1,L_SIZE), to_sfixed(0.2638,1,L_SIZE), to_sfixed(0.8359,1,L_SIZE), to_sfixed(0.6500,1,L_SIZE), to_sfixed(0.8148,1,L_SIZE), to_sfixed(0.7603,1,L_SIZE), to_sfixed(0.5394,1,L_SIZE), to_sfixed(0.7576,1,L_SIZE), to_sfixed(0.3771,1,L_SIZE), to_sfixed(0.4154,1,L_SIZE), to_sfixed(0.7310,1,L_SIZE), to_sfixed(0.7500,1,L_SIZE), to_sfixed(0.7351,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9110,1,L_SIZE), to_sfixed(0.3103,1,L_SIZE), to_sfixed(0.8204,1,L_SIZE), to_sfixed(0.6333,1,L_SIZE), to_sfixed(0.6790,1,L_SIZE), to_sfixed(0.6057,1,L_SIZE), to_sfixed(0.4980,1,L_SIZE), to_sfixed(0.4394,1,L_SIZE), to_sfixed(0.4302,1,L_SIZE), to_sfixed(0.3231,1,L_SIZE), to_sfixed(0.6433,1,L_SIZE), to_sfixed(0.7175,1,L_SIZE), to_sfixed(0.6518,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9090,1,L_SIZE), to_sfixed(0.3121,1,L_SIZE), to_sfixed(0.7461,1,L_SIZE), to_sfixed(0.6833,1,L_SIZE), to_sfixed(0.6173,1,L_SIZE), to_sfixed(0.6959,1,L_SIZE), to_sfixed(0.5866,1,L_SIZE), to_sfixed(0.3939,1,L_SIZE), to_sfixed(0.5196,1,L_SIZE), to_sfixed(0.3923,1,L_SIZE), to_sfixed(0.6082,1,L_SIZE), to_sfixed(0.8675,1,L_SIZE), to_sfixed(0.5476,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8955,1,L_SIZE), to_sfixed(0.2828,1,L_SIZE), to_sfixed(0.8793,1,L_SIZE), to_sfixed(0.5167,1,L_SIZE), to_sfixed(0.6790,1,L_SIZE), to_sfixed(0.6701,1,L_SIZE), to_sfixed(0.5276,1,L_SIZE), to_sfixed(0.5152,1,L_SIZE), to_sfixed(0.3799,1,L_SIZE), to_sfixed(0.3538,1,L_SIZE), to_sfixed(0.6374,1,L_SIZE), to_sfixed(0.6950,1,L_SIZE), to_sfixed(0.5238,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8800,1,L_SIZE), to_sfixed(0.2845,1,L_SIZE), to_sfixed(0.7895,1,L_SIZE), to_sfixed(0.6000,1,L_SIZE), to_sfixed(0.6049,1,L_SIZE), to_sfixed(0.6314,1,L_SIZE), to_sfixed(0.4783,1,L_SIZE), to_sfixed(0.4394,1,L_SIZE), to_sfixed(0.4022,1,L_SIZE), to_sfixed(0.3269,1,L_SIZE), to_sfixed(0.6550,1,L_SIZE), to_sfixed(0.6275,1,L_SIZE), to_sfixed(0.6577,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8813,1,L_SIZE), to_sfixed(0.2586,1,L_SIZE), to_sfixed(0.6502,1,L_SIZE), to_sfixed(0.5167,1,L_SIZE), to_sfixed(0.6049,1,L_SIZE), to_sfixed(0.6186,1,L_SIZE), to_sfixed(0.5197,1,L_SIZE), to_sfixed(0.4242,1,L_SIZE), to_sfixed(0.3827,1,L_SIZE), to_sfixed(0.2846,1,L_SIZE), to_sfixed(0.6901,1,L_SIZE), to_sfixed(0.6725,1,L_SIZE), to_sfixed(0.6071,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9589,1,L_SIZE), to_sfixed(0.6879,1,L_SIZE), to_sfixed(0.7771,1,L_SIZE), to_sfixed(0.4400,1,L_SIZE), to_sfixed(0.7901,1,L_SIZE), to_sfixed(0.7732,1,L_SIZE), to_sfixed(0.5984,1,L_SIZE), to_sfixed(0.3030,1,L_SIZE), to_sfixed(0.5810,1,L_SIZE), to_sfixed(0.3923,1,L_SIZE), to_sfixed(0.5205,1,L_SIZE), to_sfixed(0.8825,1,L_SIZE), to_sfixed(0.4524,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9144,1,L_SIZE), to_sfixed(0.2948,1,L_SIZE), to_sfixed(0.7152,1,L_SIZE), to_sfixed(0.5400,1,L_SIZE), to_sfixed(0.7222,1,L_SIZE), to_sfixed(0.8119,1,L_SIZE), to_sfixed(0.6476,1,L_SIZE), to_sfixed(0.5152,1,L_SIZE), to_sfixed(0.6536,1,L_SIZE), to_sfixed(0.4715,1,L_SIZE), to_sfixed(0.5556,1,L_SIZE), to_sfixed(0.8450,1,L_SIZE), to_sfixed(0.4732,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9042,1,L_SIZE), to_sfixed(0.6621,1,L_SIZE), to_sfixed(0.6563,1,L_SIZE), to_sfixed(0.6267,1,L_SIZE), to_sfixed(0.5556,1,L_SIZE), to_sfixed(0.6314,1,L_SIZE), to_sfixed(0.5276,1,L_SIZE), to_sfixed(0.4091,1,L_SIZE), to_sfixed(0.4134,1,L_SIZE), to_sfixed(0.3292,1,L_SIZE), to_sfixed(0.5322,1,L_SIZE), to_sfixed(0.7500,1,L_SIZE), to_sfixed(0.6161,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9359,1,L_SIZE), to_sfixed(0.3259,1,L_SIZE), to_sfixed(0.8019,1,L_SIZE), to_sfixed(0.5000,1,L_SIZE), to_sfixed(0.6235,1,L_SIZE), to_sfixed(0.8376,1,L_SIZE), to_sfixed(0.7008,1,L_SIZE), to_sfixed(0.2576,1,L_SIZE), to_sfixed(0.4749,1,L_SIZE), to_sfixed(0.4177,1,L_SIZE), to_sfixed(0.5146,1,L_SIZE), to_sfixed(0.8900,1,L_SIZE), to_sfixed(0.6518,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8928,1,L_SIZE), to_sfixed(0.6862,1,L_SIZE), to_sfixed(0.7090,1,L_SIZE), to_sfixed(0.5833,1,L_SIZE), to_sfixed(0.6358,1,L_SIZE), to_sfixed(0.6804,1,L_SIZE), to_sfixed(0.5177,1,L_SIZE), to_sfixed(0.4848,1,L_SIZE), to_sfixed(0.4637,1,L_SIZE), to_sfixed(0.3354,1,L_SIZE), to_sfixed(0.4795,1,L_SIZE), to_sfixed(0.7500,1,L_SIZE), to_sfixed(0.4048,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8800,1,L_SIZE), to_sfixed(0.3052,1,L_SIZE), to_sfixed(0.6502,1,L_SIZE), to_sfixed(0.5667,1,L_SIZE), to_sfixed(0.6605,1,L_SIZE), to_sfixed(0.7732,1,L_SIZE), to_sfixed(0.5906,1,L_SIZE), to_sfixed(0.4242,1,L_SIZE), to_sfixed(0.5670,1,L_SIZE), to_sfixed(0.3877,1,L_SIZE), to_sfixed(0.5146,1,L_SIZE), to_sfixed(0.8375,1,L_SIZE), to_sfixed(0.5268,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9582,1,L_SIZE), to_sfixed(0.6966,1,L_SIZE), to_sfixed(0.7554,1,L_SIZE), to_sfixed(0.6300,1,L_SIZE), to_sfixed(0.6852,1,L_SIZE), to_sfixed(0.7345,1,L_SIZE), to_sfixed(0.5217,1,L_SIZE), to_sfixed(0.4545,1,L_SIZE), to_sfixed(0.3492,1,L_SIZE), to_sfixed(0.4031,1,L_SIZE), to_sfixed(0.5088,1,L_SIZE), to_sfixed(0.8325,1,L_SIZE), to_sfixed(0.6429,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9697,1,L_SIZE), to_sfixed(0.6190,1,L_SIZE), to_sfixed(0.7059,1,L_SIZE), to_sfixed(0.5333,1,L_SIZE), to_sfixed(0.6296,1,L_SIZE), to_sfixed(0.8376,1,L_SIZE), to_sfixed(0.6240,1,L_SIZE), to_sfixed(0.4091,1,L_SIZE), to_sfixed(0.6117,1,L_SIZE), to_sfixed(0.3769,1,L_SIZE), to_sfixed(0.6082,1,L_SIZE), to_sfixed(0.8600,1,L_SIZE), to_sfixed(0.6339,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9373,1,L_SIZE), to_sfixed(0.2897,1,L_SIZE), to_sfixed(0.6563,1,L_SIZE), to_sfixed(0.5333,1,L_SIZE), to_sfixed(0.6235,1,L_SIZE), to_sfixed(0.7990,1,L_SIZE), to_sfixed(0.6673,1,L_SIZE), to_sfixed(0.3182,1,L_SIZE), to_sfixed(0.5978,1,L_SIZE), to_sfixed(0.4692,1,L_SIZE), to_sfixed(0.5322,1,L_SIZE), to_sfixed(0.8325,1,L_SIZE), to_sfixed(0.5863,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9508,1,L_SIZE), to_sfixed(0.3483,1,L_SIZE), to_sfixed(0.7430,1,L_SIZE), to_sfixed(0.6267,1,L_SIZE), to_sfixed(0.6358,1,L_SIZE), to_sfixed(0.7088,1,L_SIZE), to_sfixed(0.5748,1,L_SIZE), to_sfixed(0.4848,1,L_SIZE), to_sfixed(0.6648,1,L_SIZE), to_sfixed(0.4769,1,L_SIZE), to_sfixed(0.6257,1,L_SIZE), to_sfixed(0.6875,1,L_SIZE), to_sfixed(0.6310,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9400,1,L_SIZE), to_sfixed(0.2983,1,L_SIZE), to_sfixed(0.7028,1,L_SIZE), to_sfixed(0.5800,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(0.7423,1,L_SIZE), to_sfixed(0.6969,1,L_SIZE), to_sfixed(0.4848,1,L_SIZE), to_sfixed(0.5810,1,L_SIZE), to_sfixed(0.6846,1,L_SIZE), to_sfixed(0.6550,1,L_SIZE), to_sfixed(0.7750,1,L_SIZE), to_sfixed(0.7500,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8800,1,L_SIZE), to_sfixed(0.2983,1,L_SIZE), to_sfixed(0.6316,1,L_SIZE), to_sfixed(0.4133,1,L_SIZE), to_sfixed(0.5679,1,L_SIZE), to_sfixed(0.7010,1,L_SIZE), to_sfixed(0.6437,1,L_SIZE), to_sfixed(0.2576,1,L_SIZE), to_sfixed(0.8128,1,L_SIZE), to_sfixed(0.5538,1,L_SIZE), to_sfixed(0.6550,1,L_SIZE), to_sfixed(0.7275,1,L_SIZE), to_sfixed(0.6845,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9326,1,L_SIZE), to_sfixed(0.2845,1,L_SIZE), to_sfixed(0.8050,1,L_SIZE), to_sfixed(0.5733,1,L_SIZE), to_sfixed(0.5802,1,L_SIZE), to_sfixed(0.6314,1,L_SIZE), to_sfixed(0.5886,1,L_SIZE), to_sfixed(0.3333,1,L_SIZE), to_sfixed(0.6397,1,L_SIZE), to_sfixed(0.4308,1,L_SIZE), to_sfixed(0.7251,1,L_SIZE), to_sfixed(0.8425,1,L_SIZE), to_sfixed(0.7530,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9319,1,L_SIZE), to_sfixed(0.3017,1,L_SIZE), to_sfixed(0.7492,1,L_SIZE), to_sfixed(0.4667,1,L_SIZE), to_sfixed(0.6852,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.7362,1,L_SIZE), to_sfixed(0.4848,1,L_SIZE), to_sfixed(0.5223,1,L_SIZE), to_sfixed(0.5423,1,L_SIZE), to_sfixed(0.5906,1,L_SIZE), to_sfixed(0.8150,1,L_SIZE), to_sfixed(0.7083,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9285,1,L_SIZE), to_sfixed(0.3276,1,L_SIZE), to_sfixed(0.8297,1,L_SIZE), to_sfixed(0.5700,1,L_SIZE), to_sfixed(0.7099,1,L_SIZE), to_sfixed(0.7732,1,L_SIZE), to_sfixed(0.5492,1,L_SIZE), to_sfixed(0.5909,1,L_SIZE), to_sfixed(0.4693,1,L_SIZE), to_sfixed(0.4846,1,L_SIZE), to_sfixed(0.6608,1,L_SIZE), to_sfixed(0.7325,1,L_SIZE), to_sfixed(0.8185,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9265,1,L_SIZE), to_sfixed(0.2879,1,L_SIZE), to_sfixed(0.6966,1,L_SIZE), to_sfixed(0.5467,1,L_SIZE), to_sfixed(0.7284,1,L_SIZE), to_sfixed(0.6701,1,L_SIZE), to_sfixed(0.5709,1,L_SIZE), to_sfixed(0.3182,1,L_SIZE), to_sfixed(0.4525,1,L_SIZE), to_sfixed(0.4500,1,L_SIZE), to_sfixed(0.5380,1,L_SIZE), to_sfixed(0.8000,1,L_SIZE), to_sfixed(0.6310,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9144,1,L_SIZE), to_sfixed(0.2983,1,L_SIZE), to_sfixed(0.7616,1,L_SIZE), to_sfixed(0.6833,1,L_SIZE), to_sfixed(0.7160,1,L_SIZE), to_sfixed(0.7629,1,L_SIZE), to_sfixed(0.5472,1,L_SIZE), to_sfixed(0.3030,1,L_SIZE), to_sfixed(0.6844,1,L_SIZE), to_sfixed(0.4808,1,L_SIZE), to_sfixed(0.5731,1,L_SIZE), to_sfixed(0.7575,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9589,1,L_SIZE), to_sfixed(0.2931,1,L_SIZE), to_sfixed(0.7121,1,L_SIZE), to_sfixed(0.5433,1,L_SIZE), to_sfixed(0.7284,1,L_SIZE), to_sfixed(0.8247,1,L_SIZE), to_sfixed(0.5906,1,L_SIZE), to_sfixed(0.3939,1,L_SIZE), to_sfixed(0.5670,1,L_SIZE), to_sfixed(0.4908,1,L_SIZE), to_sfixed(0.5497,1,L_SIZE), to_sfixed(0.8275,1,L_SIZE), to_sfixed(0.5774,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8962,1,L_SIZE), to_sfixed(0.3397,1,L_SIZE), to_sfixed(0.8297,1,L_SIZE), to_sfixed(0.5600,1,L_SIZE), to_sfixed(0.6296,1,L_SIZE), to_sfixed(0.7732,1,L_SIZE), to_sfixed(0.6358,1,L_SIZE), to_sfixed(0.4697,1,L_SIZE), to_sfixed(0.4637,1,L_SIZE), to_sfixed(0.4615,1,L_SIZE), to_sfixed(0.6257,1,L_SIZE), to_sfixed(0.7100,1,L_SIZE), to_sfixed(0.7560,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9252,1,L_SIZE), to_sfixed(0.2466,1,L_SIZE), to_sfixed(0.7740,1,L_SIZE), to_sfixed(0.5567,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(0.8763,1,L_SIZE), to_sfixed(0.7224,1,L_SIZE), to_sfixed(0.2879,1,L_SIZE), to_sfixed(0.5698,1,L_SIZE), to_sfixed(0.5231,1,L_SIZE), to_sfixed(0.5205,1,L_SIZE), to_sfixed(0.7175,1,L_SIZE), to_sfixed(0.7649,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8341,1,L_SIZE), to_sfixed(0.1621,1,L_SIZE), to_sfixed(0.4211,1,L_SIZE), to_sfixed(0.3533,1,L_SIZE), to_sfixed(0.5432,1,L_SIZE), to_sfixed(0.5103,1,L_SIZE), to_sfixed(0.1122,1,L_SIZE), to_sfixed(0.4242,1,L_SIZE), to_sfixed(0.1173,1,L_SIZE), to_sfixed(0.1500,1,L_SIZE), to_sfixed(0.6140,1,L_SIZE), to_sfixed(0.4550,1,L_SIZE), to_sfixed(0.3095,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8314,1,L_SIZE), to_sfixed(0.1897,1,L_SIZE), to_sfixed(0.7059,1,L_SIZE), to_sfixed(0.5333,1,L_SIZE), to_sfixed(0.6235,1,L_SIZE), to_sfixed(0.5284,1,L_SIZE), to_sfixed(0.2146,1,L_SIZE), to_sfixed(0.9545,1,L_SIZE), to_sfixed(0.1145,1,L_SIZE), to_sfixed(0.2515,1,L_SIZE), to_sfixed(0.7310,1,L_SIZE), to_sfixed(0.4175,1,L_SIZE), to_sfixed(0.4048,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8523,1,L_SIZE), to_sfixed(0.2345,1,L_SIZE), to_sfixed(0.6254,1,L_SIZE), to_sfixed(0.5600,1,L_SIZE), to_sfixed(0.6173,1,L_SIZE), to_sfixed(0.5206,1,L_SIZE), to_sfixed(0.2776,1,L_SIZE), to_sfixed(0.8030,1,L_SIZE), to_sfixed(0.1732,1,L_SIZE), to_sfixed(0.4423,1,L_SIZE), to_sfixed(0.5731,1,L_SIZE), to_sfixed(0.3975,1,L_SIZE), to_sfixed(0.2679,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9218,1,L_SIZE), to_sfixed(0.2155,1,L_SIZE), to_sfixed(0.5944,1,L_SIZE), to_sfixed(0.6000,1,L_SIZE), to_sfixed(0.5802,1,L_SIZE), to_sfixed(0.5412,1,L_SIZE), to_sfixed(0.3524,1,L_SIZE), to_sfixed(0.4848,1,L_SIZE), to_sfixed(0.2039,1,L_SIZE), to_sfixed(0.2923,1,L_SIZE), to_sfixed(0.7193,1,L_SIZE), to_sfixed(0.6150,1,L_SIZE), to_sfixed(0.3750,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8341,1,L_SIZE), to_sfixed(0.1948,1,L_SIZE), to_sfixed(0.6687,1,L_SIZE), to_sfixed(0.6333,1,L_SIZE), to_sfixed(0.5370,1,L_SIZE), to_sfixed(0.9021,1,L_SIZE), to_sfixed(0.6102,1,L_SIZE), to_sfixed(0.2879,1,L_SIZE), to_sfixed(0.5223,1,L_SIZE), to_sfixed(0.3423,1,L_SIZE), to_sfixed(0.7135,1,L_SIZE), to_sfixed(0.7175,1,L_SIZE), to_sfixed(0.2500,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8206,1,L_SIZE), to_sfixed(0.2500,1,L_SIZE), to_sfixed(0.7833,1,L_SIZE), to_sfixed(0.6333,1,L_SIZE), to_sfixed(0.6420,1,L_SIZE), to_sfixed(0.4871,1,L_SIZE), to_sfixed(0.3445,1,L_SIZE), to_sfixed(0.6818,1,L_SIZE), to_sfixed(0.2877,1,L_SIZE), to_sfixed(0.2269,1,L_SIZE), to_sfixed(0.8480,1,L_SIZE), to_sfixed(0.5575,1,L_SIZE), to_sfixed(0.2113,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8341,1,L_SIZE), to_sfixed(0.2086,1,L_SIZE), to_sfixed(0.7926,1,L_SIZE), to_sfixed(0.6033,1,L_SIZE), to_sfixed(0.6049,1,L_SIZE), to_sfixed(0.6237,1,L_SIZE), to_sfixed(0.5217,1,L_SIZE), to_sfixed(0.5606,1,L_SIZE), to_sfixed(0.5810,1,L_SIZE), to_sfixed(0.3538,1,L_SIZE), to_sfixed(0.6959,1,L_SIZE), to_sfixed(0.5750,1,L_SIZE), to_sfixed(0.4036,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8840,1,L_SIZE), to_sfixed(0.1741,1,L_SIZE), to_sfixed(0.5263,1,L_SIZE), to_sfixed(0.5000,1,L_SIZE), to_sfixed(0.4815,1,L_SIZE), to_sfixed(0.7680,1,L_SIZE), to_sfixed(0.6260,1,L_SIZE), to_sfixed(0.3939,1,L_SIZE), to_sfixed(0.6369,1,L_SIZE), to_sfixed(0.4077,1,L_SIZE), to_sfixed(0.6550,1,L_SIZE), to_sfixed(0.7950,1,L_SIZE), to_sfixed(0.2988,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8341,1,L_SIZE), to_sfixed(0.2017,1,L_SIZE), to_sfixed(0.5944,1,L_SIZE), to_sfixed(0.6533,1,L_SIZE), to_sfixed(0.4815,1,L_SIZE), to_sfixed(0.5438,1,L_SIZE), to_sfixed(0.3937,1,L_SIZE), to_sfixed(0.4091,1,L_SIZE), to_sfixed(0.2905,1,L_SIZE), to_sfixed(0.3600,1,L_SIZE), to_sfixed(0.6550,1,L_SIZE), to_sfixed(0.8700,1,L_SIZE), to_sfixed(0.3036,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8995,1,L_SIZE), to_sfixed(0.1621,1,L_SIZE), to_sfixed(0.7307,1,L_SIZE), to_sfixed(0.5667,1,L_SIZE), to_sfixed(0.6790,1,L_SIZE), to_sfixed(0.6521,1,L_SIZE), to_sfixed(0.2559,1,L_SIZE), to_sfixed(0.8333,1,L_SIZE), to_sfixed(0.1173,1,L_SIZE), to_sfixed(0.2438,1,L_SIZE), to_sfixed(0.5965,1,L_SIZE), to_sfixed(0.4825,1,L_SIZE), to_sfixed(0.4464,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8233,1,L_SIZE), to_sfixed(0.2052,1,L_SIZE), to_sfixed(0.5418,1,L_SIZE), to_sfixed(0.5600,1,L_SIZE), to_sfixed(0.9321,1,L_SIZE), to_sfixed(0.4768,1,L_SIZE), to_sfixed(0.2520,1,L_SIZE), to_sfixed(0.2121,1,L_SIZE), to_sfixed(0.6983,1,L_SIZE), to_sfixed(0.2192,1,L_SIZE), to_sfixed(0.7485,1,L_SIZE), to_sfixed(0.7675,1,L_SIZE), to_sfixed(0.4274,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8287,1,L_SIZE), to_sfixed(0.2776,1,L_SIZE), to_sfixed(0.6842,1,L_SIZE), to_sfixed(0.6800,1,L_SIZE), to_sfixed(0.6358,1,L_SIZE), to_sfixed(0.2835,1,L_SIZE), to_sfixed(0.2008,1,L_SIZE), to_sfixed(0.5606,1,L_SIZE), to_sfixed(0.4078,1,L_SIZE), to_sfixed(0.2346,1,L_SIZE), to_sfixed(0.5298,1,L_SIZE), to_sfixed(0.4550,1,L_SIZE), to_sfixed(0.5179,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9346,1,L_SIZE), to_sfixed(0.2603,1,L_SIZE), to_sfixed(0.8266,1,L_SIZE), to_sfixed(0.8333,1,L_SIZE), to_sfixed(0.5309,1,L_SIZE), to_sfixed(0.7603,1,L_SIZE), to_sfixed(0.5630,1,L_SIZE), to_sfixed(0.3182,1,L_SIZE), to_sfixed(0.5223,1,L_SIZE), to_sfixed(0.2600,1,L_SIZE), to_sfixed(0.7953,1,L_SIZE), to_sfixed(0.7900,1,L_SIZE), to_sfixed(0.2440,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.9096,1,L_SIZE), to_sfixed(0.2862,1,L_SIZE), to_sfixed(0.6935,1,L_SIZE), to_sfixed(0.8000,1,L_SIZE), to_sfixed(0.5370,1,L_SIZE), to_sfixed(0.4845,1,L_SIZE), to_sfixed(0.3622,1,L_SIZE), to_sfixed(0.4091,1,L_SIZE), to_sfixed(0.2877,1,L_SIZE), to_sfixed(0.2877,1,L_SIZE), to_sfixed(0.5731,1,L_SIZE), to_sfixed(0.6950,1,L_SIZE), to_sfixed(0.2810,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8759,1,L_SIZE), to_sfixed(0.2879,1,L_SIZE), to_sfixed(0.8050,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.8580,1,L_SIZE), to_sfixed(0.8505,1,L_SIZE), to_sfixed(0.5689,1,L_SIZE), to_sfixed(0.3182,1,L_SIZE), to_sfixed(0.5475,1,L_SIZE), to_sfixed(0.2577,1,L_SIZE), to_sfixed(0.7661,1,L_SIZE), to_sfixed(0.8750,1,L_SIZE), to_sfixed(0.5863,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8065,1,L_SIZE), to_sfixed(0.1879,1,L_SIZE), to_sfixed(0.7121,1,L_SIZE), to_sfixed(0.7000,1,L_SIZE), to_sfixed(0.6235,1,L_SIZE), to_sfixed(0.8711,1,L_SIZE), to_sfixed(0.4213,1,L_SIZE), to_sfixed(0.1970,1,L_SIZE), to_sfixed(0.4609,1,L_SIZE), to_sfixed(0.2469,1,L_SIZE), to_sfixed(0.5789,1,L_SIZE), to_sfixed(0.7825,1,L_SIZE), to_sfixed(0.5274,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.7862,1,L_SIZE), to_sfixed(0.3241,1,L_SIZE), to_sfixed(0.5944,1,L_SIZE), to_sfixed(0.5333,1,L_SIZE), to_sfixed(0.5988,1,L_SIZE), to_sfixed(0.4149,1,L_SIZE), to_sfixed(0.3091,1,L_SIZE), to_sfixed(0.5152,1,L_SIZE), to_sfixed(0.3212,1,L_SIZE), to_sfixed(0.2923,1,L_SIZE), to_sfixed(0.7193,1,L_SIZE), to_sfixed(0.5350,1,L_SIZE), to_sfixed(0.2548,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8786,1,L_SIZE), to_sfixed(0.1552,1,L_SIZE), to_sfixed(0.5294,1,L_SIZE), to_sfixed(0.5333,1,L_SIZE), to_sfixed(0.5309,1,L_SIZE), to_sfixed(0.5026,1,L_SIZE), to_sfixed(0.3996,1,L_SIZE), to_sfixed(0.3636,1,L_SIZE), to_sfixed(0.4078,1,L_SIZE), to_sfixed(0.3538,1,L_SIZE), to_sfixed(0.6959,1,L_SIZE), to_sfixed(0.6200,1,L_SIZE), to_sfixed(0.2333,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.7984,1,L_SIZE), to_sfixed(0.4983,1,L_SIZE), to_sfixed(0.6904,1,L_SIZE), to_sfixed(0.6000,1,L_SIZE), to_sfixed(0.6914,1,L_SIZE), to_sfixed(0.4433,1,L_SIZE), to_sfixed(0.2598,1,L_SIZE), to_sfixed(0.6515,1,L_SIZE), to_sfixed(0.2654,1,L_SIZE), to_sfixed(0.2038,1,L_SIZE), to_sfixed(0.5614,1,L_SIZE), to_sfixed(0.6300,1,L_SIZE), to_sfixed(0.2976,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8314,1,L_SIZE), to_sfixed(0.1707,1,L_SIZE), to_sfixed(0.6037,1,L_SIZE), to_sfixed(0.4933,1,L_SIZE), to_sfixed(0.8395,1,L_SIZE), to_sfixed(0.4897,1,L_SIZE), to_sfixed(0.3642,1,L_SIZE), to_sfixed(0.5303,1,L_SIZE), to_sfixed(0.7709,1,L_SIZE), to_sfixed(0.2615,1,L_SIZE), to_sfixed(0.6199,1,L_SIZE), to_sfixed(0.5775,1,L_SIZE), to_sfixed(0.4464,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8564,1,L_SIZE), to_sfixed(0.6672,1,L_SIZE), to_sfixed(0.7430,1,L_SIZE), to_sfixed(0.7667,1,L_SIZE), to_sfixed(0.6235,1,L_SIZE), to_sfixed(0.7294,1,L_SIZE), to_sfixed(0.5020,1,L_SIZE), to_sfixed(0.6515,1,L_SIZE), to_sfixed(0.5447,1,L_SIZE), to_sfixed(0.1977,1,L_SIZE), to_sfixed(0.6959,1,L_SIZE), to_sfixed(0.7825,1,L_SIZE), to_sfixed(0.2756,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8092,1,L_SIZE), to_sfixed(0.1586,1,L_SIZE), to_sfixed(0.6192,1,L_SIZE), to_sfixed(0.6333,1,L_SIZE), to_sfixed(0.5309,1,L_SIZE), to_sfixed(0.6237,1,L_SIZE), to_sfixed(0.4449,1,L_SIZE), to_sfixed(0.4545,1,L_SIZE), to_sfixed(0.3994,1,L_SIZE), to_sfixed(0.1923,1,L_SIZE), to_sfixed(0.8070,1,L_SIZE), to_sfixed(0.7800,1,L_SIZE), to_sfixed(0.1655,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8577,1,L_SIZE), to_sfixed(0.3121,1,L_SIZE), to_sfixed(0.6811,1,L_SIZE), to_sfixed(0.6267,1,L_SIZE), to_sfixed(0.5309,1,L_SIZE), to_sfixed(0.5670,1,L_SIZE), to_sfixed(0.4980,1,L_SIZE), to_sfixed(0.3939,1,L_SIZE), to_sfixed(0.4944,1,L_SIZE), to_sfixed(0.3000,1,L_SIZE), to_sfixed(0.6784,1,L_SIZE), to_sfixed(0.7850,1,L_SIZE), to_sfixed(0.4250,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8146,1,L_SIZE), to_sfixed(0.1948,1,L_SIZE), to_sfixed(0.7771,1,L_SIZE), to_sfixed(0.8000,1,L_SIZE), to_sfixed(0.4815,1,L_SIZE), to_sfixed(0.5155,1,L_SIZE), to_sfixed(0.3110,1,L_SIZE), to_sfixed(0.6061,1,L_SIZE), to_sfixed(0.3911,1,L_SIZE), to_sfixed(0.1692,1,L_SIZE), to_sfixed(0.7661,1,L_SIZE), to_sfixed(0.6800,1,L_SIZE), to_sfixed(0.3750,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8800,1,L_SIZE), to_sfixed(0.6655,1,L_SIZE), to_sfixed(0.7183,1,L_SIZE), to_sfixed(0.7500,1,L_SIZE), to_sfixed(0.5247,1,L_SIZE), to_sfixed(0.4253,1,L_SIZE), to_sfixed(0.3130,1,L_SIZE), to_sfixed(0.9242,1,L_SIZE), to_sfixed(0.4525,1,L_SIZE), to_sfixed(0.3692,1,L_SIZE), to_sfixed(0.4912,1,L_SIZE), to_sfixed(0.5025,1,L_SIZE), to_sfixed(0.3065,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.7984,1,L_SIZE), to_sfixed(0.1534,1,L_SIZE), to_sfixed(0.7988,1,L_SIZE), to_sfixed(0.6000,1,L_SIZE), to_sfixed(0.5802,1,L_SIZE), to_sfixed(0.5670,1,L_SIZE), to_sfixed(0.4350,1,L_SIZE), to_sfixed(0.3333,1,L_SIZE), to_sfixed(0.6564,1,L_SIZE), to_sfixed(0.2346,1,L_SIZE), to_sfixed(0.4620,1,L_SIZE), to_sfixed(0.7700,1,L_SIZE), to_sfixed(0.3095,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8543,1,L_SIZE), to_sfixed(0.1690,1,L_SIZE), to_sfixed(0.6935,1,L_SIZE), to_sfixed(0.6000,1,L_SIZE), to_sfixed(0.6111,1,L_SIZE), to_sfixed(0.5670,1,L_SIZE), to_sfixed(0.3819,1,L_SIZE), to_sfixed(0.4545,1,L_SIZE), to_sfixed(0.4078,1,L_SIZE), to_sfixed(0.2015,1,L_SIZE), to_sfixed(0.7193,1,L_SIZE), to_sfixed(0.7900,1,L_SIZE), to_sfixed(0.2679,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8200,1,L_SIZE), to_sfixed(0.2776,1,L_SIZE), to_sfixed(0.7152,1,L_SIZE), to_sfixed(0.7600,1,L_SIZE), to_sfixed(0.5556,1,L_SIZE), to_sfixed(0.4588,1,L_SIZE), to_sfixed(0.3327,1,L_SIZE), to_sfixed(0.6515,1,L_SIZE), to_sfixed(0.4358,1,L_SIZE), to_sfixed(0.1885,1,L_SIZE), to_sfixed(0.7778,1,L_SIZE), to_sfixed(0.5650,1,L_SIZE), to_sfixed(0.2946,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.7856,1,L_SIZE), to_sfixed(0.2879,1,L_SIZE), to_sfixed(0.8111,1,L_SIZE), to_sfixed(0.8667,1,L_SIZE), to_sfixed(0.5432,1,L_SIZE), to_sfixed(0.4948,1,L_SIZE), to_sfixed(0.3169,1,L_SIZE), to_sfixed(0.6061,1,L_SIZE), to_sfixed(0.3743,1,L_SIZE), to_sfixed(0.2000,1,L_SIZE), to_sfixed(0.7953,1,L_SIZE), to_sfixed(0.8025,1,L_SIZE), to_sfixed(0.3345,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.7849,1,L_SIZE), to_sfixed(0.3552,1,L_SIZE), to_sfixed(0.7616,1,L_SIZE), to_sfixed(0.7200,1,L_SIZE), to_sfixed(0.5185,1,L_SIZE), to_sfixed(0.5026,1,L_SIZE), to_sfixed(0.3327,1,L_SIZE), to_sfixed(0.7273,1,L_SIZE), to_sfixed(0.3771,1,L_SIZE), to_sfixed(0.2154,1,L_SIZE), to_sfixed(0.5848,1,L_SIZE), to_sfixed(0.6875,1,L_SIZE), to_sfixed(0.4048,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8146,1,L_SIZE), to_sfixed(0.2293,1,L_SIZE), to_sfixed(0.7121,1,L_SIZE), to_sfixed(0.7867,1,L_SIZE), to_sfixed(0.4321,1,L_SIZE), to_sfixed(0.5670,1,L_SIZE), to_sfixed(0.3130,1,L_SIZE), to_sfixed(0.6364,1,L_SIZE), to_sfixed(0.3855,1,L_SIZE), to_sfixed(0.1338,1,L_SIZE), to_sfixed(0.6257,1,L_SIZE), to_sfixed(0.8025,1,L_SIZE), to_sfixed(0.3720,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8146,1,L_SIZE), to_sfixed(0.3155,1,L_SIZE), to_sfixed(0.7183,1,L_SIZE), to_sfixed(0.6167,1,L_SIZE), to_sfixed(0.5000,1,L_SIZE), to_sfixed(0.4124,1,L_SIZE), to_sfixed(0.2953,1,L_SIZE), to_sfixed(0.7879,1,L_SIZE), to_sfixed(0.4581,1,L_SIZE), to_sfixed(0.1846,1,L_SIZE), to_sfixed(0.6316,1,L_SIZE), to_sfixed(0.5675,1,L_SIZE), to_sfixed(0.2857,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8092,1,L_SIZE), to_sfixed(0.2603,1,L_SIZE), to_sfixed(0.7492,1,L_SIZE), to_sfixed(0.7333,1,L_SIZE), to_sfixed(0.5309,1,L_SIZE), to_sfixed(0.3737,1,L_SIZE), to_sfixed(0.2461,1,L_SIZE), to_sfixed(0.7576,1,L_SIZE), to_sfixed(0.4553,1,L_SIZE), to_sfixed(0.2769,1,L_SIZE), to_sfixed(0.6140,1,L_SIZE), to_sfixed(0.6625,1,L_SIZE), to_sfixed(0.2679,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8557,1,L_SIZE), to_sfixed(0.2638,1,L_SIZE), to_sfixed(0.6997,1,L_SIZE), to_sfixed(0.6900,1,L_SIZE), to_sfixed(0.4938,1,L_SIZE), to_sfixed(0.3557,1,L_SIZE), to_sfixed(0.2874,1,L_SIZE), to_sfixed(0.8788,1,L_SIZE), to_sfixed(0.4525,1,L_SIZE), to_sfixed(0.2346,1,L_SIZE), to_sfixed(0.5614,1,L_SIZE), to_sfixed(0.5150,1,L_SIZE), to_sfixed(0.2946,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8287,1,L_SIZE), to_sfixed(0.4879,1,L_SIZE), to_sfixed(0.6873,1,L_SIZE), to_sfixed(0.6000,1,L_SIZE), to_sfixed(0.5432,1,L_SIZE), to_sfixed(0.6314,1,L_SIZE), to_sfixed(0.4429,1,L_SIZE), to_sfixed(0.3788,1,L_SIZE), to_sfixed(0.5559,1,L_SIZE), to_sfixed(0.1654,1,L_SIZE), to_sfixed(0.6725,1,L_SIZE), to_sfixed(0.8250,1,L_SIZE), to_sfixed(0.1726,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.7835,1,L_SIZE), to_sfixed(0.3431,1,L_SIZE), to_sfixed(0.7059,1,L_SIZE), to_sfixed(0.6000,1,L_SIZE), to_sfixed(0.6049,1,L_SIZE), to_sfixed(0.7784,1,L_SIZE), to_sfixed(0.4449,1,L_SIZE), to_sfixed(0.2576,1,L_SIZE), to_sfixed(0.3771,1,L_SIZE), to_sfixed(0.2500,1,L_SIZE), to_sfixed(0.6784,1,L_SIZE), to_sfixed(0.7400,1,L_SIZE), to_sfixed(0.2054,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8409,1,L_SIZE), to_sfixed(0.2621,1,L_SIZE), to_sfixed(0.6811,1,L_SIZE), to_sfixed(0.6333,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.6443,1,L_SIZE), to_sfixed(0.4469,1,L_SIZE), to_sfixed(0.4848,1,L_SIZE), to_sfixed(0.9162,1,L_SIZE), to_sfixed(0.2000,1,L_SIZE), to_sfixed(0.6784,1,L_SIZE), to_sfixed(0.6575,1,L_SIZE), to_sfixed(0.5577,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.7964,1,L_SIZE), to_sfixed(0.3655,1,L_SIZE), to_sfixed(0.8483,1,L_SIZE), to_sfixed(0.7167,1,L_SIZE), to_sfixed(0.8272,1,L_SIZE), to_sfixed(0.4124,1,L_SIZE), to_sfixed(0.1949,1,L_SIZE), to_sfixed(0.2121,1,L_SIZE), to_sfixed(0.4358,1,L_SIZE), to_sfixed(0.1923,1,L_SIZE), to_sfixed(0.5556,1,L_SIZE), to_sfixed(0.5650,1,L_SIZE), to_sfixed(0.3720,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8287,1,L_SIZE), to_sfixed(0.2431,1,L_SIZE), to_sfixed(0.6130,1,L_SIZE), to_sfixed(0.5333,1,L_SIZE), to_sfixed(0.5247,1,L_SIZE), to_sfixed(0.6572,1,L_SIZE), to_sfixed(0.4921,1,L_SIZE), to_sfixed(0.4394,1,L_SIZE), to_sfixed(0.4944,1,L_SIZE), to_sfixed(0.2231,1,L_SIZE), to_sfixed(0.7193,1,L_SIZE), to_sfixed(0.6850,1,L_SIZE), to_sfixed(0.2548,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8341,1,L_SIZE), to_sfixed(0.1845,1,L_SIZE), to_sfixed(0.6502,1,L_SIZE), to_sfixed(0.6167,1,L_SIZE), to_sfixed(0.5432,1,L_SIZE), to_sfixed(0.9072,1,L_SIZE), to_sfixed(0.7382,1,L_SIZE), to_sfixed(0.3636,1,L_SIZE), to_sfixed(0.5447,1,L_SIZE), to_sfixed(0.3462,1,L_SIZE), to_sfixed(0.6082,1,L_SIZE), to_sfixed(0.6925,1,L_SIZE), to_sfixed(0.3929,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8287,1,L_SIZE), to_sfixed(0.5466,1,L_SIZE), to_sfixed(0.6842,1,L_SIZE), to_sfixed(0.6000,1,L_SIZE), to_sfixed(0.5432,1,L_SIZE), to_sfixed(0.7345,1,L_SIZE), to_sfixed(0.5886,1,L_SIZE), to_sfixed(0.6818,1,L_SIZE), to_sfixed(0.7849,1,L_SIZE), to_sfixed(0.1769,1,L_SIZE), to_sfixed(0.8304,1,L_SIZE), to_sfixed(0.7075,1,L_SIZE), to_sfixed(0.2417,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8146,1,L_SIZE), to_sfixed(0.3586,1,L_SIZE), to_sfixed(0.5263,1,L_SIZE), to_sfixed(0.5833,1,L_SIZE), to_sfixed(0.5988,1,L_SIZE), to_sfixed(0.5747,1,L_SIZE), to_sfixed(0.4272,1,L_SIZE), to_sfixed(0.3939,1,L_SIZE), to_sfixed(0.3911,1,L_SIZE), to_sfixed(0.2538,1,L_SIZE), to_sfixed(0.7427,1,L_SIZE), to_sfixed(0.7400,1,L_SIZE), to_sfixed(0.4226,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8496,1,L_SIZE), to_sfixed(0.2310,1,L_SIZE), to_sfixed(0.5882,1,L_SIZE), to_sfixed(0.6167,1,L_SIZE), to_sfixed(0.5432,1,L_SIZE), to_sfixed(0.3737,1,L_SIZE), to_sfixed(0.2677,1,L_SIZE), to_sfixed(0.4394,1,L_SIZE), to_sfixed(0.3771,1,L_SIZE), to_sfixed(0.1885,1,L_SIZE), to_sfixed(0.6082,1,L_SIZE), to_sfixed(0.6925,1,L_SIZE), to_sfixed(0.3345,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8321,1,L_SIZE), to_sfixed(0.4224,1,L_SIZE), to_sfixed(0.7616,1,L_SIZE), to_sfixed(0.7000,1,L_SIZE), to_sfixed(0.6049,1,L_SIZE), to_sfixed(0.6598,1,L_SIZE), to_sfixed(0.4154,1,L_SIZE), to_sfixed(0.5152,1,L_SIZE), to_sfixed(0.3659,1,L_SIZE), to_sfixed(0.2154,1,L_SIZE), to_sfixed(0.4678,1,L_SIZE), to_sfixed(0.8450,1,L_SIZE), to_sfixed(0.2607,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.7970,1,L_SIZE), to_sfixed(0.2966,1,L_SIZE), to_sfixed(0.5820,1,L_SIZE), to_sfixed(0.6500,1,L_SIZE), to_sfixed(0.5309,1,L_SIZE), to_sfixed(0.6443,1,L_SIZE), to_sfixed(0.3228,1,L_SIZE), to_sfixed(0.5606,1,L_SIZE), to_sfixed(0.3966,1,L_SIZE), to_sfixed(0.1585,1,L_SIZE), to_sfixed(0.5497,1,L_SIZE), to_sfixed(0.6100,1,L_SIZE), to_sfixed(0.2470,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8436,1,L_SIZE), to_sfixed(0.2983,1,L_SIZE), to_sfixed(0.6130,1,L_SIZE), to_sfixed(0.6833,1,L_SIZE), to_sfixed(0.5247,1,L_SIZE), to_sfixed(0.5670,1,L_SIZE), to_sfixed(0.3780,1,L_SIZE), to_sfixed(0.4848,1,L_SIZE), to_sfixed(0.4134,1,L_SIZE), to_sfixed(0.2262,1,L_SIZE), to_sfixed(0.6082,1,L_SIZE), to_sfixed(0.8925,1,L_SIZE), to_sfixed(0.4000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8375,1,L_SIZE), to_sfixed(0.4397,1,L_SIZE), to_sfixed(0.7028,1,L_SIZE), to_sfixed(0.7333,1,L_SIZE), to_sfixed(0.5556,1,L_SIZE), to_sfixed(0.4330,1,L_SIZE), to_sfixed(0.3622,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.3966,1,L_SIZE), to_sfixed(0.2077,1,L_SIZE), to_sfixed(0.5029,1,L_SIZE), to_sfixed(0.8250,1,L_SIZE), to_sfixed(0.1875,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8260,1,L_SIZE), to_sfixed(0.2983,1,L_SIZE), to_sfixed(0.6563,1,L_SIZE), to_sfixed(0.6333,1,L_SIZE), to_sfixed(0.4938,1,L_SIZE), to_sfixed(0.4253,1,L_SIZE), to_sfixed(0.3996,1,L_SIZE), to_sfixed(0.5606,1,L_SIZE), to_sfixed(0.4553,1,L_SIZE), to_sfixed(0.2615,1,L_SIZE), to_sfixed(0.5848,1,L_SIZE), to_sfixed(0.7925,1,L_SIZE), to_sfixed(0.3036,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8577,1,L_SIZE), to_sfixed(0.3017,1,L_SIZE), to_sfixed(0.7059,1,L_SIZE), to_sfixed(0.7500,1,L_SIZE), to_sfixed(0.5185,1,L_SIZE), to_sfixed(0.3557,1,L_SIZE), to_sfixed(0.3465,1,L_SIZE), to_sfixed(0.7273,1,L_SIZE), to_sfixed(0.4553,1,L_SIZE), to_sfixed(0.2538,1,L_SIZE), to_sfixed(0.5146,1,L_SIZE), to_sfixed(0.6050,1,L_SIZE), to_sfixed(0.2905,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8240,1,L_SIZE), to_sfixed(0.2224,1,L_SIZE), to_sfixed(0.6006,1,L_SIZE), to_sfixed(0.6333,1,L_SIZE), to_sfixed(0.5679,1,L_SIZE), to_sfixed(0.6082,1,L_SIZE), to_sfixed(0.4016,1,L_SIZE), to_sfixed(0.5909,1,L_SIZE), to_sfixed(0.5810,1,L_SIZE), to_sfixed(0.2077,1,L_SIZE), to_sfixed(0.5029,1,L_SIZE), to_sfixed(0.7550,1,L_SIZE), to_sfixed(0.1857,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.7829,1,L_SIZE), to_sfixed(0.2328,1,L_SIZE), to_sfixed(0.8359,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(0.5802,1,L_SIZE), to_sfixed(0.7062,1,L_SIZE), to_sfixed(0.5748,1,L_SIZE), to_sfixed(0.4394,1,L_SIZE), to_sfixed(0.6955,1,L_SIZE), to_sfixed(0.2038,1,L_SIZE), to_sfixed(0.5614,1,L_SIZE), to_sfixed(0.8150,1,L_SIZE), to_sfixed(0.4048,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.7728,1,L_SIZE), to_sfixed(0.6448,1,L_SIZE), to_sfixed(0.5635,1,L_SIZE), to_sfixed(0.6500,1,L_SIZE), to_sfixed(0.6605,1,L_SIZE), to_sfixed(0.8196,1,L_SIZE), to_sfixed(0.5079,1,L_SIZE), to_sfixed(0.3636,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.2231,1,L_SIZE), to_sfixed(0.4386,1,L_SIZE), to_sfixed(0.7025,1,L_SIZE), to_sfixed(0.3345,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8442,1,L_SIZE), to_sfixed(0.4190,1,L_SIZE), to_sfixed(0.6718,1,L_SIZE), to_sfixed(0.7000,1,L_SIZE), to_sfixed(0.5432,1,L_SIZE), to_sfixed(0.6572,1,L_SIZE), to_sfixed(0.4469,1,L_SIZE), to_sfixed(0.3939,1,L_SIZE), to_sfixed(0.3408,1,L_SIZE), to_sfixed(0.1538,1,L_SIZE), to_sfixed(0.5263,1,L_SIZE), to_sfixed(0.6950,1,L_SIZE), to_sfixed(0.1935,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.7930,1,L_SIZE), to_sfixed(0.4621,1,L_SIZE), to_sfixed(0.9040,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(0.6358,1,L_SIZE), to_sfixed(0.4510,1,L_SIZE), to_sfixed(0.3996,1,L_SIZE), to_sfixed(0.9091,1,L_SIZE), to_sfixed(0.2933,1,L_SIZE), to_sfixed(0.2923,1,L_SIZE), to_sfixed(0.7193,1,L_SIZE), to_sfixed(0.6250,1,L_SIZE), to_sfixed(0.3613,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.7694,1,L_SIZE), to_sfixed(0.1276,1,L_SIZE), to_sfixed(0.7740,1,L_SIZE), to_sfixed(0.7000,1,L_SIZE), to_sfixed(0.5432,1,L_SIZE), to_sfixed(0.6392,1,L_SIZE), to_sfixed(0.3957,1,L_SIZE), to_sfixed(0.6364,1,L_SIZE), to_sfixed(0.4022,1,L_SIZE), to_sfixed(0.2369,1,L_SIZE), to_sfixed(0.6433,1,L_SIZE), to_sfixed(0.5775,1,L_SIZE), to_sfixed(0.2583,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8146,1,L_SIZE), to_sfixed(0.2397,1,L_SIZE), to_sfixed(0.7740,1,L_SIZE), to_sfixed(0.7500,1,L_SIZE), to_sfixed(0.5185,1,L_SIZE), to_sfixed(0.6598,1,L_SIZE), to_sfixed(0.4508,1,L_SIZE), to_sfixed(0.6515,1,L_SIZE), to_sfixed(0.2905,1,L_SIZE), to_sfixed(0.2231,1,L_SIZE), to_sfixed(0.5439,1,L_SIZE), to_sfixed(0.7975,1,L_SIZE), to_sfixed(0.2292,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.7438,1,L_SIZE), to_sfixed(0.2603,1,L_SIZE), to_sfixed(0.6811,1,L_SIZE), to_sfixed(0.7167,1,L_SIZE), to_sfixed(0.5247,1,L_SIZE), to_sfixed(0.6340,1,L_SIZE), to_sfixed(0.4272,1,L_SIZE), to_sfixed(0.7879,1,L_SIZE), to_sfixed(0.5615,1,L_SIZE), to_sfixed(0.1462,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.7175,1,L_SIZE), to_sfixed(0.2423,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.7970,1,L_SIZE), to_sfixed(0.2534,1,L_SIZE), to_sfixed(0.6161,1,L_SIZE), to_sfixed(0.6933,1,L_SIZE), to_sfixed(0.5309,1,L_SIZE), to_sfixed(0.5103,1,L_SIZE), to_sfixed(0.3150,1,L_SIZE), to_sfixed(0.4545,1,L_SIZE), to_sfixed(0.4274,1,L_SIZE), to_sfixed(0.1500,1,L_SIZE), to_sfixed(0.5556,1,L_SIZE), to_sfixed(0.8325,1,L_SIZE), to_sfixed(0.2946,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8375,1,L_SIZE), to_sfixed(0.2776,1,L_SIZE), to_sfixed(0.6780,1,L_SIZE), to_sfixed(0.7500,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(0.5155,1,L_SIZE), to_sfixed(0.4114,1,L_SIZE), to_sfixed(0.5152,1,L_SIZE), to_sfixed(0.4497,1,L_SIZE), to_sfixed(0.1585,1,L_SIZE), to_sfixed(0.6199,1,L_SIZE), to_sfixed(0.7400,1,L_SIZE), to_sfixed(0.2054,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8611,1,L_SIZE), to_sfixed(0.5914,1,L_SIZE), to_sfixed(0.6130,1,L_SIZE), to_sfixed(0.5333,1,L_SIZE), to_sfixed(0.4938,1,L_SIZE), to_sfixed(0.4201,1,L_SIZE), to_sfixed(0.2461,1,L_SIZE), to_sfixed(0.6515,1,L_SIZE), to_sfixed(0.2318,1,L_SIZE), to_sfixed(0.2615,1,L_SIZE), to_sfixed(0.4094,1,L_SIZE), to_sfixed(0.5300,1,L_SIZE), to_sfixed(0.2214,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8092,1,L_SIZE), to_sfixed(0.5914,1,L_SIZE), to_sfixed(0.6192,1,L_SIZE), to_sfixed(0.6333,1,L_SIZE), to_sfixed(0.5370,1,L_SIZE), to_sfixed(0.5155,1,L_SIZE), to_sfixed(0.3228,1,L_SIZE), to_sfixed(0.5606,1,L_SIZE), to_sfixed(0.5223,1,L_SIZE), to_sfixed(0.0985,1,L_SIZE), to_sfixed(0.5439,1,L_SIZE), to_sfixed(0.7625,1,L_SIZE), to_sfixed(0.3357,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.7721,1,L_SIZE), to_sfixed(0.4138,1,L_SIZE), to_sfixed(0.7492,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(0.5926,1,L_SIZE), to_sfixed(0.7474,1,L_SIZE), to_sfixed(0.5492,1,L_SIZE), to_sfixed(0.4848,1,L_SIZE), to_sfixed(0.5112,1,L_SIZE), to_sfixed(0.2500,1,L_SIZE), to_sfixed(0.4678,1,L_SIZE), to_sfixed(0.8475,1,L_SIZE), to_sfixed(0.3720,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.7795,1,L_SIZE), to_sfixed(0.3534,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.9500,1,L_SIZE), to_sfixed(0.7346,1,L_SIZE), to_sfixed(0.8196,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.7121,1,L_SIZE), to_sfixed(0.5223,1,L_SIZE), to_sfixed(0.4615,1,L_SIZE), to_sfixed(0.5439,1,L_SIZE), to_sfixed(0.9225,1,L_SIZE), to_sfixed(0.2768,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8375,1,L_SIZE), to_sfixed(0.7638,1,L_SIZE), to_sfixed(0.8452,1,L_SIZE), to_sfixed(0.8833,1,L_SIZE), to_sfixed(0.6296,1,L_SIZE), to_sfixed(0.5670,1,L_SIZE), to_sfixed(0.4193,1,L_SIZE), to_sfixed(0.6515,1,L_SIZE), to_sfixed(0.4777,1,L_SIZE), to_sfixed(0.1600,1,L_SIZE), to_sfixed(0.5380,1,L_SIZE), to_sfixed(0.7800,1,L_SIZE), to_sfixed(0.2173,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8800,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.6594,1,L_SIZE), to_sfixed(0.7167,1,L_SIZE), to_sfixed(0.5309,1,L_SIZE), to_sfixed(0.6753,1,L_SIZE), to_sfixed(0.5217,1,L_SIZE), to_sfixed(0.4545,1,L_SIZE), to_sfixed(0.5615,1,L_SIZE), to_sfixed(0.2000,1,L_SIZE), to_sfixed(0.4269,1,L_SIZE), to_sfixed(0.7750,1,L_SIZE), to_sfixed(0.2262,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8004,1,L_SIZE), to_sfixed(0.7431,1,L_SIZE), to_sfixed(0.7399,1,L_SIZE), to_sfixed(0.7000,1,L_SIZE), to_sfixed(0.5062,1,L_SIZE), to_sfixed(0.7371,1,L_SIZE), to_sfixed(0.5965,1,L_SIZE), to_sfixed(0.3182,1,L_SIZE), to_sfixed(0.8128,1,L_SIZE), to_sfixed(0.2154,1,L_SIZE), to_sfixed(0.4386,1,L_SIZE), to_sfixed(0.9100,1,L_SIZE), to_sfixed(0.2262,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8139,1,L_SIZE), to_sfixed(0.3724,1,L_SIZE), to_sfixed(0.6718,1,L_SIZE), to_sfixed(0.7000,1,L_SIZE), to_sfixed(0.5247,1,L_SIZE), to_sfixed(0.6701,1,L_SIZE), to_sfixed(0.5217,1,L_SIZE), to_sfixed(0.5606,1,L_SIZE), to_sfixed(0.3771,1,L_SIZE), to_sfixed(0.2123,1,L_SIZE), to_sfixed(0.5029,1,L_SIZE), to_sfixed(0.8200,1,L_SIZE), to_sfixed(0.2250,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8382,1,L_SIZE), to_sfixed(0.2638,1,L_SIZE), to_sfixed(0.7090,1,L_SIZE), to_sfixed(0.7167,1,L_SIZE), to_sfixed(0.5309,1,L_SIZE), to_sfixed(0.7062,1,L_SIZE), to_sfixed(0.6201,1,L_SIZE), to_sfixed(0.5909,1,L_SIZE), to_sfixed(0.4944,1,L_SIZE), to_sfixed(0.3031,1,L_SIZE), to_sfixed(0.4035,1,L_SIZE), to_sfixed(0.7100,1,L_SIZE), to_sfixed(0.2095,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.7950,1,L_SIZE), to_sfixed(0.3672,1,L_SIZE), to_sfixed(0.8607,1,L_SIZE), to_sfixed(0.9500,1,L_SIZE), to_sfixed(0.5679,1,L_SIZE), to_sfixed(0.5490,1,L_SIZE), to_sfixed(0.4409,1,L_SIZE), to_sfixed(0.8788,1,L_SIZE), to_sfixed(0.4916,1,L_SIZE), to_sfixed(0.2308,1,L_SIZE), to_sfixed(0.5673,1,L_SIZE), to_sfixed(0.6100,1,L_SIZE), to_sfixed(0.2774,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8341,1,L_SIZE), to_sfixed(0.2810,1,L_SIZE), to_sfixed(0.7121,1,L_SIZE), to_sfixed(0.8167,1,L_SIZE), to_sfixed(0.5432,1,L_SIZE), to_sfixed(0.5722,1,L_SIZE), to_sfixed(0.4823,1,L_SIZE), to_sfixed(0.6061,1,L_SIZE), to_sfixed(0.5307,1,L_SIZE), to_sfixed(0.1631,1,L_SIZE), to_sfixed(0.5205,1,L_SIZE), to_sfixed(0.6950,1,L_SIZE), to_sfixed(0.2036,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8119,1,L_SIZE), to_sfixed(0.7414,1,L_SIZE), to_sfixed(0.7368,1,L_SIZE), to_sfixed(0.7333,1,L_SIZE), to_sfixed(0.4938,1,L_SIZE), to_sfixed(0.5412,1,L_SIZE), to_sfixed(0.3445,1,L_SIZE), to_sfixed(0.6364,1,L_SIZE), to_sfixed(0.3771,1,L_SIZE), to_sfixed(0.2000,1,L_SIZE), to_sfixed(0.4620,1,L_SIZE), to_sfixed(0.6425,1,L_SIZE), to_sfixed(0.3452,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE)),
					(to_sfixed(0.8672,1,L_SIZE), to_sfixed(0.2328,1,L_SIZE), to_sfixed(0.7183,1,L_SIZE), to_sfixed(0.6000,1,L_SIZE), to_sfixed(0.7531,1,L_SIZE), to_sfixed(0.3892,1,L_SIZE), to_sfixed(0.2461,1,L_SIZE), to_sfixed(0.3182,1,L_SIZE), to_sfixed(0.2626,1,L_SIZE), to_sfixed(0.3154,1,L_SIZE), to_sfixed(0.4444,1,L_SIZE), to_sfixed(0.3225,1,L_SIZE), to_sfixed(0.3750,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8685,1,L_SIZE), to_sfixed(0.5155,1,L_SIZE), to_sfixed(0.7430,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(0.6420,1,L_SIZE), to_sfixed(0.3351,1,L_SIZE), to_sfixed(0.2402,1,L_SIZE), to_sfixed(0.3636,1,L_SIZE), to_sfixed(0.2318,1,L_SIZE), to_sfixed(0.4154,1,L_SIZE), to_sfixed(0.4327,1,L_SIZE), to_sfixed(0.3550,1,L_SIZE), to_sfixed(0.3155,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8638,1,L_SIZE), to_sfixed(0.3983,1,L_SIZE), to_sfixed(0.7430,1,L_SIZE), to_sfixed(0.8000,1,L_SIZE), to_sfixed(0.6049,1,L_SIZE), to_sfixed(0.2964,1,L_SIZE), to_sfixed(0.2146,1,L_SIZE), to_sfixed(0.4091,1,L_SIZE), to_sfixed(0.2318,1,L_SIZE), to_sfixed(0.4385,1,L_SIZE), to_sfixed(0.3860,1,L_SIZE), to_sfixed(0.3400,1,L_SIZE), to_sfixed(0.3333,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8564,1,L_SIZE), to_sfixed(0.6121,1,L_SIZE), to_sfixed(0.7307,1,L_SIZE), to_sfixed(0.7167,1,L_SIZE), to_sfixed(0.6543,1,L_SIZE), to_sfixed(0.4381,1,L_SIZE), to_sfixed(0.2362,1,L_SIZE), to_sfixed(0.2576,1,L_SIZE), to_sfixed(0.2346,1,L_SIZE), to_sfixed(0.3846,1,L_SIZE), to_sfixed(0.4561,1,L_SIZE), to_sfixed(0.3225,1,L_SIZE), to_sfixed(0.3571,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8436,1,L_SIZE), to_sfixed(0.2138,1,L_SIZE), to_sfixed(0.6966,1,L_SIZE), to_sfixed(0.5833,1,L_SIZE), to_sfixed(0.5247,1,L_SIZE), to_sfixed(0.5155,1,L_SIZE), to_sfixed(0.1142,1,L_SIZE), to_sfixed(0.9091,1,L_SIZE), to_sfixed(0.3492,1,L_SIZE), to_sfixed(0.4192,1,L_SIZE), to_sfixed(0.4386,1,L_SIZE), to_sfixed(0.3775,1,L_SIZE), to_sfixed(0.3869,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8496,1,L_SIZE), to_sfixed(0.4241,1,L_SIZE), to_sfixed(0.6811,1,L_SIZE), to_sfixed(0.6167,1,L_SIZE), to_sfixed(0.5802,1,L_SIZE), to_sfixed(0.4175,1,L_SIZE), to_sfixed(0.1299,1,L_SIZE), to_sfixed(0.9545,1,L_SIZE), to_sfixed(0.2626,1,L_SIZE), to_sfixed(0.5462,1,L_SIZE), to_sfixed(0.4269,1,L_SIZE), to_sfixed(0.3950,1,L_SIZE), to_sfixed(0.4137,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8260,1,L_SIZE), to_sfixed(0.8138,1,L_SIZE), to_sfixed(0.7864,1,L_SIZE), to_sfixed(0.7000,1,L_SIZE), to_sfixed(0.5494,1,L_SIZE), to_sfixed(0.3557,1,L_SIZE), to_sfixed(0.0925,1,L_SIZE), to_sfixed(0.8030,1,L_SIZE), to_sfixed(0.2235,1,L_SIZE), to_sfixed(0.2962,1,L_SIZE), to_sfixed(0.4386,1,L_SIZE), to_sfixed(0.3175,1,L_SIZE), to_sfixed(0.4286,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8449,1,L_SIZE), to_sfixed(0.9500,1,L_SIZE), to_sfixed(0.8173,1,L_SIZE), to_sfixed(0.8333,1,L_SIZE), to_sfixed(0.5926,1,L_SIZE), to_sfixed(0.4613,1,L_SIZE), to_sfixed(0.1181,1,L_SIZE), to_sfixed(0.9545,1,L_SIZE), to_sfixed(0.3073,1,L_SIZE), to_sfixed(0.3846,1,L_SIZE), to_sfixed(0.4795,1,L_SIZE), to_sfixed(0.4225,1,L_SIZE), to_sfixed(0.3065,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.9096,1,L_SIZE), to_sfixed(0.6190,1,L_SIZE), to_sfixed(0.6780,1,L_SIZE), to_sfixed(0.6500,1,L_SIZE), to_sfixed(0.5432,1,L_SIZE), to_sfixed(0.4175,1,L_SIZE), to_sfixed(0.0945,1,L_SIZE), to_sfixed(0.8788,1,L_SIZE), to_sfixed(0.2458,1,L_SIZE), to_sfixed(0.4385,1,L_SIZE), to_sfixed(0.4737,1,L_SIZE), to_sfixed(0.4550,1,L_SIZE), to_sfixed(0.3452,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8658,1,L_SIZE), to_sfixed(0.5103,1,L_SIZE), to_sfixed(0.8080,1,L_SIZE), to_sfixed(0.8000,1,L_SIZE), to_sfixed(0.6235,1,L_SIZE), to_sfixed(0.5979,1,L_SIZE), to_sfixed(0.1181,1,L_SIZE), to_sfixed(0.8030,1,L_SIZE), to_sfixed(0.2263,1,L_SIZE), to_sfixed(0.3785,1,L_SIZE), to_sfixed(0.5205,1,L_SIZE), to_sfixed(0.5375,1,L_SIZE), to_sfixed(0.3512,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8719,1,L_SIZE), to_sfixed(0.4845,1,L_SIZE), to_sfixed(0.8359,1,L_SIZE), to_sfixed(0.7000,1,L_SIZE), to_sfixed(0.5926,1,L_SIZE), to_sfixed(0.3969,1,L_SIZE), to_sfixed(0.0984,1,L_SIZE), to_sfixed(0.8030,1,L_SIZE), to_sfixed(0.2095,1,L_SIZE), to_sfixed(0.3538,1,L_SIZE), to_sfixed(0.4503,1,L_SIZE), to_sfixed(0.5775,1,L_SIZE), to_sfixed(0.3571,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.9009,1,L_SIZE), to_sfixed(0.4414,1,L_SIZE), to_sfixed(0.7276,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(0.5494,1,L_SIZE), to_sfixed(0.3608,1,L_SIZE), to_sfixed(0.0984,1,L_SIZE), to_sfixed(0.5606,1,L_SIZE), to_sfixed(0.1788,1,L_SIZE), to_sfixed(0.4308,1,L_SIZE), to_sfixed(0.4094,1,L_SIZE), to_sfixed(0.6175,1,L_SIZE), to_sfixed(0.4643,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.9117,1,L_SIZE), to_sfixed(0.5466,1,L_SIZE), to_sfixed(0.8421,1,L_SIZE), to_sfixed(0.7833,1,L_SIZE), to_sfixed(0.5988,1,L_SIZE), to_sfixed(0.3995,1,L_SIZE), to_sfixed(0.1024,1,L_SIZE), to_sfixed(0.7576,1,L_SIZE), to_sfixed(0.1536,1,L_SIZE), to_sfixed(0.3346,1,L_SIZE), to_sfixed(0.5205,1,L_SIZE), to_sfixed(0.5150,1,L_SIZE), to_sfixed(0.3095,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.9184,1,L_SIZE), to_sfixed(0.8534,1,L_SIZE), to_sfixed(0.7276,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(0.5679,1,L_SIZE), to_sfixed(0.5155,1,L_SIZE), to_sfixed(0.1575,1,L_SIZE), to_sfixed(0.7121,1,L_SIZE), to_sfixed(0.2849,1,L_SIZE), to_sfixed(0.3385,1,L_SIZE), to_sfixed(0.5322,1,L_SIZE), to_sfixed(0.5125,1,L_SIZE), to_sfixed(0.3274,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8260,1,L_SIZE), to_sfixed(0.6690,1,L_SIZE), to_sfixed(0.6811,1,L_SIZE), to_sfixed(0.6167,1,L_SIZE), to_sfixed(0.6914,1,L_SIZE), to_sfixed(0.3557,1,L_SIZE), to_sfixed(0.1535,1,L_SIZE), to_sfixed(0.4394,1,L_SIZE), to_sfixed(0.3184,1,L_SIZE), to_sfixed(0.6315,1,L_SIZE), to_sfixed(0.3801,1,L_SIZE), to_sfixed(0.5000,1,L_SIZE), to_sfixed(0.5089,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8874,1,L_SIZE), to_sfixed(0.6155,1,L_SIZE), to_sfixed(0.6656,1,L_SIZE), to_sfixed(0.7000,1,L_SIZE), to_sfixed(0.6296,1,L_SIZE), to_sfixed(0.3866,1,L_SIZE), to_sfixed(0.1083,1,L_SIZE), to_sfixed(0.6515,1,L_SIZE), to_sfixed(0.3631,1,L_SIZE), to_sfixed(0.3077,1,L_SIZE), to_sfixed(0.3509,1,L_SIZE), to_sfixed(0.4200,1,L_SIZE), to_sfixed(0.4940,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.9359,1,L_SIZE), to_sfixed(0.8690,1,L_SIZE), to_sfixed(0.6904,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(0.4938,1,L_SIZE), to_sfixed(0.2526,1,L_SIZE), to_sfixed(0.0669,1,L_SIZE), to_sfixed(0.6061,1,L_SIZE), to_sfixed(0.1899,1,L_SIZE), to_sfixed(0.3769,1,L_SIZE), to_sfixed(0.3392,1,L_SIZE), to_sfixed(0.3325,1,L_SIZE), to_sfixed(0.2470,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8678,1,L_SIZE), to_sfixed(0.7948,1,L_SIZE), to_sfixed(0.7678,1,L_SIZE), to_sfixed(0.7167,1,L_SIZE), to_sfixed(0.5309,1,L_SIZE), to_sfixed(0.4381,1,L_SIZE), to_sfixed(0.1280,1,L_SIZE), to_sfixed(0.7121,1,L_SIZE), to_sfixed(0.2402,1,L_SIZE), to_sfixed(0.5885,1,L_SIZE), to_sfixed(0.3158,1,L_SIZE), to_sfixed(0.4650,1,L_SIZE), to_sfixed(0.3720,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8982,1,L_SIZE), to_sfixed(0.5586,1,L_SIZE), to_sfixed(0.7368,1,L_SIZE), to_sfixed(0.7167,1,L_SIZE), to_sfixed(0.5679,1,L_SIZE), to_sfixed(0.4974,1,L_SIZE), to_sfixed(0.1496,1,L_SIZE), to_sfixed(0.6818,1,L_SIZE), to_sfixed(0.3492,1,L_SIZE), to_sfixed(0.6477,1,L_SIZE), to_sfixed(0.3216,1,L_SIZE), to_sfixed(0.4050,1,L_SIZE), to_sfixed(0.3869,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8820,1,L_SIZE), to_sfixed(0.6724,1,L_SIZE), to_sfixed(0.7307,1,L_SIZE), to_sfixed(0.7167,1,L_SIZE), to_sfixed(0.6975,1,L_SIZE), to_sfixed(0.3634,1,L_SIZE), to_sfixed(0.2736,1,L_SIZE), to_sfixed(0.5152,1,L_SIZE), to_sfixed(0.3184,1,L_SIZE), to_sfixed(0.7231,1,L_SIZE), to_sfixed(0.3333,1,L_SIZE), to_sfixed(0.3325,1,L_SIZE), to_sfixed(0.3274,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.9103,1,L_SIZE), to_sfixed(0.5379,1,L_SIZE), to_sfixed(0.8111,1,L_SIZE), to_sfixed(0.8000,1,L_SIZE), to_sfixed(0.7593,1,L_SIZE), to_sfixed(0.3608,1,L_SIZE), to_sfixed(0.3091,1,L_SIZE), to_sfixed(0.3333,1,L_SIZE), to_sfixed(0.3492,1,L_SIZE), to_sfixed(0.6615,1,L_SIZE), to_sfixed(0.3450,1,L_SIZE), to_sfixed(0.3250,1,L_SIZE), to_sfixed(0.2976,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8624,1,L_SIZE), to_sfixed(0.4603,1,L_SIZE), to_sfixed(0.7678,1,L_SIZE), to_sfixed(0.7333,1,L_SIZE), to_sfixed(0.6914,1,L_SIZE), to_sfixed(0.3814,1,L_SIZE), to_sfixed(0.2677,1,L_SIZE), to_sfixed(0.3636,1,L_SIZE), to_sfixed(0.3520,1,L_SIZE), to_sfixed(0.8308,1,L_SIZE), to_sfixed(0.2807,1,L_SIZE), to_sfixed(0.3675,1,L_SIZE), to_sfixed(0.2857,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8840,1,L_SIZE), to_sfixed(0.3276,1,L_SIZE), to_sfixed(0.8514,1,L_SIZE), to_sfixed(0.8500,1,L_SIZE), to_sfixed(0.7160,1,L_SIZE), to_sfixed(0.5670,1,L_SIZE), to_sfixed(0.2520,1,L_SIZE), to_sfixed(0.3939,1,L_SIZE), to_sfixed(0.4358,1,L_SIZE), to_sfixed(0.5462,1,L_SIZE), to_sfixed(0.3567,1,L_SIZE), to_sfixed(0.3325,1,L_SIZE), to_sfixed(0.2530,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8921,1,L_SIZE), to_sfixed(0.5690,1,L_SIZE), to_sfixed(0.7059,1,L_SIZE), to_sfixed(0.6167,1,L_SIZE), to_sfixed(0.6049,1,L_SIZE), to_sfixed(0.4639,1,L_SIZE), to_sfixed(0.1634,1,L_SIZE), to_sfixed(0.9242,1,L_SIZE), to_sfixed(0.5223,1,L_SIZE), to_sfixed(0.8092,1,L_SIZE), to_sfixed(0.3275,1,L_SIZE), to_sfixed(0.3775,1,L_SIZE), to_sfixed(0.4018,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8483,1,L_SIZE), to_sfixed(0.2224,1,L_SIZE), to_sfixed(0.6502,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(0.6358,1,L_SIZE), to_sfixed(0.3814,1,L_SIZE), to_sfixed(0.1142,1,L_SIZE), to_sfixed(0.8030,1,L_SIZE), to_sfixed(0.3911,1,L_SIZE), to_sfixed(0.5846,1,L_SIZE), to_sfixed(0.3392,1,L_SIZE), to_sfixed(0.3875,1,L_SIZE), to_sfixed(0.3810,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8881,1,L_SIZE), to_sfixed(0.8948,1,L_SIZE), to_sfixed(0.7183,1,L_SIZE), to_sfixed(0.7333,1,L_SIZE), to_sfixed(0.5741,1,L_SIZE), to_sfixed(0.4485,1,L_SIZE), to_sfixed(0.1240,1,L_SIZE), to_sfixed(0.9242,1,L_SIZE), to_sfixed(0.4330,1,L_SIZE), to_sfixed(0.6077,1,L_SIZE), to_sfixed(0.3509,1,L_SIZE), to_sfixed(0.3700,1,L_SIZE), to_sfixed(0.4315,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.9332,1,L_SIZE), to_sfixed(0.7103,1,L_SIZE), to_sfixed(0.7368,1,L_SIZE), to_sfixed(0.6500,1,L_SIZE), to_sfixed(0.5494,1,L_SIZE), to_sfixed(0.4639,1,L_SIZE), to_sfixed(0.1634,1,L_SIZE), to_sfixed(0.7273,1,L_SIZE), to_sfixed(0.4358,1,L_SIZE), to_sfixed(0.6931,1,L_SIZE), to_sfixed(0.3333,1,L_SIZE), to_sfixed(0.4100,1,L_SIZE), to_sfixed(0.2857,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8395,1,L_SIZE), to_sfixed(0.5224,1,L_SIZE), to_sfixed(0.8173,1,L_SIZE), to_sfixed(0.9000,1,L_SIZE), to_sfixed(0.5988,1,L_SIZE), to_sfixed(0.4897,1,L_SIZE), to_sfixed(0.1142,1,L_SIZE), to_sfixed(0.9545,1,L_SIZE), to_sfixed(0.3184,1,L_SIZE), to_sfixed(0.5769,1,L_SIZE), to_sfixed(0.3918,1,L_SIZE), to_sfixed(0.4325,1,L_SIZE), to_sfixed(0.5238,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.9670,1,L_SIZE), to_sfixed(0.2897,1,L_SIZE), to_sfixed(0.8359,1,L_SIZE), to_sfixed(0.8333,1,L_SIZE), to_sfixed(0.6049,1,L_SIZE), to_sfixed(0.7216,1,L_SIZE), to_sfixed(0.2579,1,L_SIZE), to_sfixed(0.8030,1,L_SIZE), to_sfixed(0.7542,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE), to_sfixed(0.3333,1,L_SIZE), to_sfixed(0.4900,1,L_SIZE), to_sfixed(0.3929,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.9090,1,L_SIZE), to_sfixed(0.2879,1,L_SIZE), to_sfixed(0.8173,1,L_SIZE), to_sfixed(0.7500,1,L_SIZE), to_sfixed(0.5494,1,L_SIZE), to_sfixed(0.6701,1,L_SIZE), to_sfixed(0.2165,1,L_SIZE), to_sfixed(0.7879,1,L_SIZE), to_sfixed(0.6397,1,L_SIZE), to_sfixed(0.9038,1,L_SIZE), to_sfixed(0.3333,1,L_SIZE), to_sfixed(0.4450,1,L_SIZE), to_sfixed(0.3690,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8334,1,L_SIZE), to_sfixed(0.6603,1,L_SIZE), to_sfixed(0.7368,1,L_SIZE), to_sfixed(0.7000,1,L_SIZE), to_sfixed(0.5432,1,L_SIZE), to_sfixed(0.5928,1,L_SIZE), to_sfixed(0.1811,1,L_SIZE), to_sfixed(0.7576,1,L_SIZE), to_sfixed(0.2905,1,L_SIZE), to_sfixed(0.5885,1,L_SIZE), to_sfixed(0.3275,1,L_SIZE), to_sfixed(0.3950,1,L_SIZE), to_sfixed(0.3095,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.9231,1,L_SIZE), to_sfixed(0.5621,1,L_SIZE), to_sfixed(0.7864,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(0.6605,1,L_SIZE), to_sfixed(0.4716,1,L_SIZE), to_sfixed(0.1102,1,L_SIZE), to_sfixed(0.7576,1,L_SIZE), to_sfixed(0.2235,1,L_SIZE), to_sfixed(0.4523,1,L_SIZE), to_sfixed(0.5614,1,L_SIZE), to_sfixed(0.4550,1,L_SIZE), to_sfixed(0.4048,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8665,1,L_SIZE), to_sfixed(0.5638,1,L_SIZE), to_sfixed(0.7988,1,L_SIZE), to_sfixed(0.7333,1,L_SIZE), to_sfixed(0.6543,1,L_SIZE), to_sfixed(0.4253,1,L_SIZE), to_sfixed(0.1181,1,L_SIZE), to_sfixed(0.9091,1,L_SIZE), to_sfixed(0.2682,1,L_SIZE), to_sfixed(0.4292,1,L_SIZE), to_sfixed(0.5088,1,L_SIZE), to_sfixed(0.5275,1,L_SIZE), to_sfixed(0.3393,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8739,1,L_SIZE), to_sfixed(0.5948,1,L_SIZE), to_sfixed(0.7276,1,L_SIZE), to_sfixed(0.6167,1,L_SIZE), to_sfixed(0.6543,1,L_SIZE), to_sfixed(0.3582,1,L_SIZE), to_sfixed(0.1378,1,L_SIZE), to_sfixed(0.6061,1,L_SIZE), to_sfixed(0.2626,1,L_SIZE), to_sfixed(0.4062,1,L_SIZE), to_sfixed(0.3977,1,L_SIZE), to_sfixed(0.4375,1,L_SIZE), to_sfixed(0.4018,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.9292,1,L_SIZE), to_sfixed(0.4759,1,L_SIZE), to_sfixed(0.7121,1,L_SIZE), to_sfixed(0.7333,1,L_SIZE), to_sfixed(0.5556,1,L_SIZE), to_sfixed(0.3479,1,L_SIZE), to_sfixed(0.1339,1,L_SIZE), to_sfixed(0.6212,1,L_SIZE), to_sfixed(0.2877,1,L_SIZE), to_sfixed(0.7369,1,L_SIZE), to_sfixed(0.4094,1,L_SIZE), to_sfixed(0.4200,1,L_SIZE), to_sfixed(0.3661,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.9258,1,L_SIZE), to_sfixed(0.7517,1,L_SIZE), to_sfixed(0.6997,1,L_SIZE), to_sfixed(0.7500,1,L_SIZE), to_sfixed(0.5432,1,L_SIZE), to_sfixed(0.3299,1,L_SIZE), to_sfixed(0.0925,1,L_SIZE), to_sfixed(0.7879,1,L_SIZE), to_sfixed(0.3212,1,L_SIZE), to_sfixed(0.5092,1,L_SIZE), to_sfixed(0.4561,1,L_SIZE), to_sfixed(0.4375,1,L_SIZE), to_sfixed(0.3095,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.9069,1,L_SIZE), to_sfixed(0.6379,1,L_SIZE), to_sfixed(0.8050,1,L_SIZE), to_sfixed(0.7667,1,L_SIZE), to_sfixed(0.6852,1,L_SIZE), to_sfixed(0.4381,1,L_SIZE), to_sfixed(0.1811,1,L_SIZE), to_sfixed(0.6515,1,L_SIZE), to_sfixed(0.4078,1,L_SIZE), to_sfixed(0.8215,1,L_SIZE), to_sfixed(0.4971,1,L_SIZE), to_sfixed(0.3900,1,L_SIZE), to_sfixed(0.4137,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8645,1,L_SIZE), to_sfixed(0.5810,1,L_SIZE), to_sfixed(0.7121,1,L_SIZE), to_sfixed(0.6500,1,L_SIZE), to_sfixed(0.5432,1,L_SIZE), to_sfixed(0.3814,1,L_SIZE), to_sfixed(0.1299,1,L_SIZE), to_sfixed(0.6061,1,L_SIZE), to_sfixed(0.2709,1,L_SIZE), to_sfixed(0.7892,1,L_SIZE), to_sfixed(0.4211,1,L_SIZE), to_sfixed(0.4375,1,L_SIZE), to_sfixed(0.4077,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.9157,1,L_SIZE), to_sfixed(0.4448,1,L_SIZE), to_sfixed(0.8328,1,L_SIZE), to_sfixed(0.8167,1,L_SIZE), to_sfixed(0.6481,1,L_SIZE), to_sfixed(0.3995,1,L_SIZE), to_sfixed(0.1654,1,L_SIZE), to_sfixed(0.5909,1,L_SIZE), to_sfixed(0.4302,1,L_SIZE), to_sfixed(0.6662,1,L_SIZE), to_sfixed(0.4327,1,L_SIZE), to_sfixed(0.4500,1,L_SIZE), to_sfixed(0.4464,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.9036,1,L_SIZE), to_sfixed(0.7931,1,L_SIZE), to_sfixed(0.8854,1,L_SIZE), to_sfixed(0.8333,1,L_SIZE), to_sfixed(0.6914,1,L_SIZE), to_sfixed(0.5103,1,L_SIZE), to_sfixed(0.1890,1,L_SIZE), to_sfixed(0.4091,1,L_SIZE), to_sfixed(0.3101,1,L_SIZE), to_sfixed(0.6538,1,L_SIZE), to_sfixed(0.3918,1,L_SIZE), to_sfixed(0.4800,1,L_SIZE), to_sfixed(0.3750,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8227,1,L_SIZE), to_sfixed(0.5224,1,L_SIZE), to_sfixed(0.7183,1,L_SIZE), to_sfixed(0.6333,1,L_SIZE), to_sfixed(0.5926,1,L_SIZE), to_sfixed(0.3222,1,L_SIZE), to_sfixed(0.0965,1,L_SIZE), to_sfixed(0.6061,1,L_SIZE), to_sfixed(0.2039,1,L_SIZE), to_sfixed(0.4231,1,L_SIZE), to_sfixed(0.3860,1,L_SIZE), to_sfixed(0.4575,1,L_SIZE), to_sfixed(0.3036,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8611,1,L_SIZE), to_sfixed(0.4121,1,L_SIZE), to_sfixed(0.7059,1,L_SIZE), to_sfixed(0.6500,1,L_SIZE), to_sfixed(0.5309,1,L_SIZE), to_sfixed(0.3582,1,L_SIZE), to_sfixed(0.1004,1,L_SIZE), to_sfixed(0.7273,1,L_SIZE), to_sfixed(0.1788,1,L_SIZE), to_sfixed(0.7615,1,L_SIZE), to_sfixed(0.3333,1,L_SIZE), to_sfixed(0.4075,1,L_SIZE), to_sfixed(0.2798,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.9548,1,L_SIZE), to_sfixed(0.4328,1,L_SIZE), to_sfixed(0.7678,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(0.5617,1,L_SIZE), to_sfixed(0.4330,1,L_SIZE), to_sfixed(0.1378,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(0.3464,1,L_SIZE), to_sfixed(0.7462,1,L_SIZE), to_sfixed(0.3626,1,L_SIZE), to_sfixed(0.4275,1,L_SIZE), to_sfixed(0.3929,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.9245,1,L_SIZE), to_sfixed(0.9741,1,L_SIZE), to_sfixed(0.7585,1,L_SIZE), to_sfixed(0.6833,1,L_SIZE), to_sfixed(0.5864,1,L_SIZE), to_sfixed(0.4330,1,L_SIZE), to_sfixed(0.1201,1,L_SIZE), to_sfixed(0.7879,1,L_SIZE), to_sfixed(0.2961,1,L_SIZE), to_sfixed(0.5923,1,L_SIZE), to_sfixed(0.3743,1,L_SIZE), to_sfixed(0.4350,1,L_SIZE), to_sfixed(0.4405,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.9036,1,L_SIZE), to_sfixed(0.6741,1,L_SIZE), to_sfixed(0.7678,1,L_SIZE), to_sfixed(0.7667,1,L_SIZE), to_sfixed(0.6296,1,L_SIZE), to_sfixed(0.4639,1,L_SIZE), to_sfixed(0.1476,1,L_SIZE), to_sfixed(0.6515,1,L_SIZE), to_sfixed(0.3939,1,L_SIZE), to_sfixed(0.5615,1,L_SIZE), to_sfixed(0.4094,1,L_SIZE), to_sfixed(0.3900,1,L_SIZE), to_sfixed(0.4464,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8948,1,L_SIZE), to_sfixed(0.7379,1,L_SIZE), to_sfixed(0.6997,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(0.7407,1,L_SIZE), to_sfixed(0.4098,1,L_SIZE), to_sfixed(0.1358,1,L_SIZE), to_sfixed(0.6515,1,L_SIZE), to_sfixed(0.3771,1,L_SIZE), to_sfixed(0.7846,1,L_SIZE), to_sfixed(0.3450,1,L_SIZE), to_sfixed(0.3900,1,L_SIZE), to_sfixed(0.4970,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.8881,1,L_SIZE), to_sfixed(0.4466,1,L_SIZE), to_sfixed(0.7337,1,L_SIZE), to_sfixed(0.6667,1,L_SIZE), to_sfixed(0.7407,1,L_SIZE), to_sfixed(0.4253,1,L_SIZE), to_sfixed(0.1339,1,L_SIZE), to_sfixed(0.8030,1,L_SIZE), to_sfixed(0.4078,1,L_SIZE), to_sfixed(0.7154,1,L_SIZE), to_sfixed(0.3509,1,L_SIZE), to_sfixed(0.4050,1,L_SIZE), to_sfixed(0.5000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE)),
					(to_sfixed(0.9528,1,L_SIZE), to_sfixed(0.7069,1,L_SIZE), to_sfixed(0.8483,1,L_SIZE), to_sfixed(0.8167,1,L_SIZE), to_sfixed(0.5926,1,L_SIZE), to_sfixed(0.5284,1,L_SIZE), to_sfixed(0.1496,1,L_SIZE), to_sfixed(0.8485,1,L_SIZE), to_sfixed(0.3771,1,L_SIZE), to_sfixed(0.7077,1,L_SIZE), to_sfixed(0.3567,1,L_SIZE), to_sfixed(0.4000,1,L_SIZE), to_sfixed(0.3333,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(0.0000,1,L_SIZE), to_sfixed(1.0000,1,L_SIZE))
				);


  -- Signals
	signal	INPUT													: ARRAY_OF_SFIXED (0 to (PERCEPTRONS_INPUT-1));
	signal	FROM_LOOKUP											: ARRAY_OF_SFIXED (0 to (PERCEPTRONS_HIDDEN-1));
	signal	OUTPUT												: ARRAY_OF_SFIXED (0 to (PERCEPTRONS_HIDDEN-1));
	  -- Signals
	signal IN_UNSIGNED						: unsigned(7 downto 0);
	signal LOOKUP_TABLE_K 					: unsigned(7 downto 0);
	signal LOOKUP_TABLE_OUT 				: INPUT_LOOKUP_ARRAY;
	signal LOOKUP_TABLE_OUT_CONSTRAINED	: INPUT_CONSTRAINED_SFIXED_ARRAY;
	signal UNIT_DELAY_OUT					: INPUT_CONSTRAINED_SFIXED_ARRAY;
	
	
--=============================================================================
-- architecture begin
--=============================================================================	
	begin
		IN_UNSIGNED <= unsigned(SAMPLE_NUMBER);
		LOOKUP_TABLE_K <= -- Make sure no index will fall out of boundary
			to_unsigned(0, 8) when IN_UNSIGNED <= 0 
		else
			to_unsigned(SAMPLE_SIZE, 8) when IN_UNSIGNED >= SAMPLE_SIZE 
		else
			IN_UNSIGNED;
  
		LOOKUP_TABLE_OUT <= INPUTS_TABLE(to_integer(LOOKUP_TABLE_K));
		
		
		GEN_PROPER_OUTPUT: 
		for I in 0 to (PERCEPTRONS_INPUT-1+PERCEPTRONS_OUTPUT) generate
			LOOKUP_TABLE_OUT_CONSTRAINED(I)<=
				resize(LOOKUP_TABLE_OUT(I),U_SIZE,L_SIZE);
								
		end generate GEN_PROPER_OUTPUT;

		UNIT_DELAY_PROCESS : process (clk)
			
			begin
				if CLK'event and CLK = '1' then
				UNIT_DELAY_OUT <= LOOKUP_TABLE_OUT_CONSTRAINED;
				end if;
		
		end process UNIT_DELAY_PROCESS;


		SELECTED_INPUT <= UNIT_DELAY_OUT;
end RTL;
--=============================================================================
-- architecture end
--=============================================================================
