--=============================================================================
--    This file is part of FPGA_NEURAL-Network.
--
--    FPGA_NEURAL-Network is free software: you can redistribute it and/or 
--    modify it under the terms of the GNU General Public License as published 
--    by the Free Software Foundation, either version 3 of the License, or
--    (at your option) any later version.
--
--    FPGA_NEURAL-Network is distributed in the hope that it will be useful,
--    but WITHOUT ANY WARRANTY; without even the implied warranty of
--    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--    GNU General Public License for more details.
--
--    You should have received a copy of the GNU General Public License
--    along with FPGA_NEURAL-Network.  
--		if not, see <http://www.gnu.org/licenses/>.

--=============================================================================
--	FILE NAME			: SIGMOID_ROM.vhd
--	PROJECT				: FPGA_NEURAL-Network
--	ENTITY				: SIGMOID_ROM
--	ARCHITECTURE		: rtl
--=============================================================================
--	AUTORS(s)			: Agostini, N;
--	DEPARTMENT      	: Electrical Engineering (UFRGS)
--	DATE					: Dec 14, 2014
--=============================================================================
--	Description:
--	
--=============================================================================

library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all; -- is the to unsigned really required????
	use work.fixed_pkg.all; -- ieee_proposed for compatibility version
	use work.NN_TYPES_pkg.all;
	use work.SIGMOID_ROM_pkg.all;

--=============================================================================
-- Entity declaration for SIGMOID_ROM
--=============================================================================
entity SIGMOID_ROM is 
	port (
		clk				:	in std_logic;
		X_VALUE 			: 	in std_logic_vector (13 downto 0);
		Y_VALUE			: 	out CONSTRAINED_SFIXED
	);
end SIGMOID_ROM;

--=============================================================================
-- architecture declaration
--=============================================================================
architecture RTL of SIGMOID_ROM is
-- Constants

			-- This constant has 16384 values
			constant TAN_SIG : TAN_SIG_VECTOR := (
				to_sfixed(-0.9951,1,L_SIZE),
				to_sfixed(-0.9951,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9950,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9949,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9948,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9947,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9946,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9945,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9944,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9943,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9942,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9941,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9940,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9939,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9938,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9937,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9936,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9935,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9934,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9933,1,L_SIZE),
				to_sfixed(-0.9932,1,L_SIZE),
				to_sfixed(-0.9932,1,L_SIZE),
				to_sfixed(-0.9932,1,L_SIZE),
				to_sfixed(-0.9932,1,L_SIZE),
				to_sfixed(-0.9932,1,L_SIZE),
				to_sfixed(-0.9932,1,L_SIZE),
				to_sfixed(-0.9932,1,L_SIZE),
				to_sfixed(-0.9932,1,L_SIZE),
				to_sfixed(-0.9932,1,L_SIZE),
				to_sfixed(-0.9932,1,L_SIZE),
				to_sfixed(-0.9932,1,L_SIZE),
				to_sfixed(-0.9932,1,L_SIZE),
				to_sfixed(-0.9932,1,L_SIZE),
				to_sfixed(-0.9932,1,L_SIZE),
				to_sfixed(-0.9932,1,L_SIZE),
				to_sfixed(-0.9932,1,L_SIZE),
				to_sfixed(-0.9932,1,L_SIZE),
				to_sfixed(-0.9932,1,L_SIZE),
				to_sfixed(-0.9932,1,L_SIZE),
				to_sfixed(-0.9932,1,L_SIZE),
				to_sfixed(-0.9931,1,L_SIZE),
				to_sfixed(-0.9931,1,L_SIZE),
				to_sfixed(-0.9931,1,L_SIZE),
				to_sfixed(-0.9931,1,L_SIZE),
				to_sfixed(-0.9931,1,L_SIZE),
				to_sfixed(-0.9931,1,L_SIZE),
				to_sfixed(-0.9931,1,L_SIZE),
				to_sfixed(-0.9931,1,L_SIZE),
				to_sfixed(-0.9931,1,L_SIZE),
				to_sfixed(-0.9931,1,L_SIZE),
				to_sfixed(-0.9931,1,L_SIZE),
				to_sfixed(-0.9931,1,L_SIZE),
				to_sfixed(-0.9931,1,L_SIZE),
				to_sfixed(-0.9931,1,L_SIZE),
				to_sfixed(-0.9931,1,L_SIZE),
				to_sfixed(-0.9931,1,L_SIZE),
				to_sfixed(-0.9931,1,L_SIZE),
				to_sfixed(-0.9931,1,L_SIZE),
				to_sfixed(-0.9931,1,L_SIZE),
				to_sfixed(-0.9931,1,L_SIZE),
				to_sfixed(-0.9930,1,L_SIZE),
				to_sfixed(-0.9930,1,L_SIZE),
				to_sfixed(-0.9930,1,L_SIZE),
				to_sfixed(-0.9930,1,L_SIZE),
				to_sfixed(-0.9930,1,L_SIZE),
				to_sfixed(-0.9930,1,L_SIZE),
				to_sfixed(-0.9930,1,L_SIZE),
				to_sfixed(-0.9930,1,L_SIZE),
				to_sfixed(-0.9930,1,L_SIZE),
				to_sfixed(-0.9930,1,L_SIZE),
				to_sfixed(-0.9930,1,L_SIZE),
				to_sfixed(-0.9930,1,L_SIZE),
				to_sfixed(-0.9930,1,L_SIZE),
				to_sfixed(-0.9930,1,L_SIZE),
				to_sfixed(-0.9930,1,L_SIZE),
				to_sfixed(-0.9930,1,L_SIZE),
				to_sfixed(-0.9930,1,L_SIZE),
				to_sfixed(-0.9930,1,L_SIZE),
				to_sfixed(-0.9930,1,L_SIZE),
				to_sfixed(-0.9929,1,L_SIZE),
				to_sfixed(-0.9929,1,L_SIZE),
				to_sfixed(-0.9929,1,L_SIZE),
				to_sfixed(-0.9929,1,L_SIZE),
				to_sfixed(-0.9929,1,L_SIZE),
				to_sfixed(-0.9929,1,L_SIZE),
				to_sfixed(-0.9929,1,L_SIZE),
				to_sfixed(-0.9929,1,L_SIZE),
				to_sfixed(-0.9929,1,L_SIZE),
				to_sfixed(-0.9929,1,L_SIZE),
				to_sfixed(-0.9929,1,L_SIZE),
				to_sfixed(-0.9929,1,L_SIZE),
				to_sfixed(-0.9929,1,L_SIZE),
				to_sfixed(-0.9929,1,L_SIZE),
				to_sfixed(-0.9929,1,L_SIZE),
				to_sfixed(-0.9929,1,L_SIZE),
				to_sfixed(-0.9929,1,L_SIZE),
				to_sfixed(-0.9929,1,L_SIZE),
				to_sfixed(-0.9929,1,L_SIZE),
				to_sfixed(-0.9928,1,L_SIZE),
				to_sfixed(-0.9928,1,L_SIZE),
				to_sfixed(-0.9928,1,L_SIZE),
				to_sfixed(-0.9928,1,L_SIZE),
				to_sfixed(-0.9928,1,L_SIZE),
				to_sfixed(-0.9928,1,L_SIZE),
				to_sfixed(-0.9928,1,L_SIZE),
				to_sfixed(-0.9928,1,L_SIZE),
				to_sfixed(-0.9928,1,L_SIZE),
				to_sfixed(-0.9928,1,L_SIZE),
				to_sfixed(-0.9928,1,L_SIZE),
				to_sfixed(-0.9928,1,L_SIZE),
				to_sfixed(-0.9928,1,L_SIZE),
				to_sfixed(-0.9928,1,L_SIZE),
				to_sfixed(-0.9928,1,L_SIZE),
				to_sfixed(-0.9928,1,L_SIZE),
				to_sfixed(-0.9928,1,L_SIZE),
				to_sfixed(-0.9928,1,L_SIZE),
				to_sfixed(-0.9928,1,L_SIZE),
				to_sfixed(-0.9927,1,L_SIZE),
				to_sfixed(-0.9927,1,L_SIZE),
				to_sfixed(-0.9927,1,L_SIZE),
				to_sfixed(-0.9927,1,L_SIZE),
				to_sfixed(-0.9927,1,L_SIZE),
				to_sfixed(-0.9927,1,L_SIZE),
				to_sfixed(-0.9927,1,L_SIZE),
				to_sfixed(-0.9927,1,L_SIZE),
				to_sfixed(-0.9927,1,L_SIZE),
				to_sfixed(-0.9927,1,L_SIZE),
				to_sfixed(-0.9927,1,L_SIZE),
				to_sfixed(-0.9927,1,L_SIZE),
				to_sfixed(-0.9927,1,L_SIZE),
				to_sfixed(-0.9927,1,L_SIZE),
				to_sfixed(-0.9927,1,L_SIZE),
				to_sfixed(-0.9927,1,L_SIZE),
				to_sfixed(-0.9927,1,L_SIZE),
				to_sfixed(-0.9927,1,L_SIZE),
				to_sfixed(-0.9927,1,L_SIZE),
				to_sfixed(-0.9926,1,L_SIZE),
				to_sfixed(-0.9926,1,L_SIZE),
				to_sfixed(-0.9926,1,L_SIZE),
				to_sfixed(-0.9926,1,L_SIZE),
				to_sfixed(-0.9926,1,L_SIZE),
				to_sfixed(-0.9926,1,L_SIZE),
				to_sfixed(-0.9926,1,L_SIZE),
				to_sfixed(-0.9926,1,L_SIZE),
				to_sfixed(-0.9926,1,L_SIZE),
				to_sfixed(-0.9926,1,L_SIZE),
				to_sfixed(-0.9926,1,L_SIZE),
				to_sfixed(-0.9926,1,L_SIZE),
				to_sfixed(-0.9926,1,L_SIZE),
				to_sfixed(-0.9926,1,L_SIZE),
				to_sfixed(-0.9926,1,L_SIZE),
				to_sfixed(-0.9926,1,L_SIZE),
				to_sfixed(-0.9926,1,L_SIZE),
				to_sfixed(-0.9926,1,L_SIZE),
				to_sfixed(-0.9926,1,L_SIZE),
				to_sfixed(-0.9925,1,L_SIZE),
				to_sfixed(-0.9925,1,L_SIZE),
				to_sfixed(-0.9925,1,L_SIZE),
				to_sfixed(-0.9925,1,L_SIZE),
				to_sfixed(-0.9925,1,L_SIZE),
				to_sfixed(-0.9925,1,L_SIZE),
				to_sfixed(-0.9925,1,L_SIZE),
				to_sfixed(-0.9925,1,L_SIZE),
				to_sfixed(-0.9925,1,L_SIZE),
				to_sfixed(-0.9925,1,L_SIZE),
				to_sfixed(-0.9925,1,L_SIZE),
				to_sfixed(-0.9925,1,L_SIZE),
				to_sfixed(-0.9925,1,L_SIZE),
				to_sfixed(-0.9925,1,L_SIZE),
				to_sfixed(-0.9925,1,L_SIZE),
				to_sfixed(-0.9925,1,L_SIZE),
				to_sfixed(-0.9925,1,L_SIZE),
				to_sfixed(-0.9925,1,L_SIZE),
				to_sfixed(-0.9924,1,L_SIZE),
				to_sfixed(-0.9924,1,L_SIZE),
				to_sfixed(-0.9924,1,L_SIZE),
				to_sfixed(-0.9924,1,L_SIZE),
				to_sfixed(-0.9924,1,L_SIZE),
				to_sfixed(-0.9924,1,L_SIZE),
				to_sfixed(-0.9924,1,L_SIZE),
				to_sfixed(-0.9924,1,L_SIZE),
				to_sfixed(-0.9924,1,L_SIZE),
				to_sfixed(-0.9924,1,L_SIZE),
				to_sfixed(-0.9924,1,L_SIZE),
				to_sfixed(-0.9924,1,L_SIZE),
				to_sfixed(-0.9924,1,L_SIZE),
				to_sfixed(-0.9924,1,L_SIZE),
				to_sfixed(-0.9924,1,L_SIZE),
				to_sfixed(-0.9924,1,L_SIZE),
				to_sfixed(-0.9924,1,L_SIZE),
				to_sfixed(-0.9924,1,L_SIZE),
				to_sfixed(-0.9923,1,L_SIZE),
				to_sfixed(-0.9923,1,L_SIZE),
				to_sfixed(-0.9923,1,L_SIZE),
				to_sfixed(-0.9923,1,L_SIZE),
				to_sfixed(-0.9923,1,L_SIZE),
				to_sfixed(-0.9923,1,L_SIZE),
				to_sfixed(-0.9923,1,L_SIZE),
				to_sfixed(-0.9923,1,L_SIZE),
				to_sfixed(-0.9923,1,L_SIZE),
				to_sfixed(-0.9923,1,L_SIZE),
				to_sfixed(-0.9923,1,L_SIZE),
				to_sfixed(-0.9923,1,L_SIZE),
				to_sfixed(-0.9923,1,L_SIZE),
				to_sfixed(-0.9923,1,L_SIZE),
				to_sfixed(-0.9923,1,L_SIZE),
				to_sfixed(-0.9923,1,L_SIZE),
				to_sfixed(-0.9923,1,L_SIZE),
				to_sfixed(-0.9923,1,L_SIZE),
				to_sfixed(-0.9922,1,L_SIZE),
				to_sfixed(-0.9922,1,L_SIZE),
				to_sfixed(-0.9922,1,L_SIZE),
				to_sfixed(-0.9922,1,L_SIZE),
				to_sfixed(-0.9922,1,L_SIZE),
				to_sfixed(-0.9922,1,L_SIZE),
				to_sfixed(-0.9922,1,L_SIZE),
				to_sfixed(-0.9922,1,L_SIZE),
				to_sfixed(-0.9922,1,L_SIZE),
				to_sfixed(-0.9922,1,L_SIZE),
				to_sfixed(-0.9922,1,L_SIZE),
				to_sfixed(-0.9922,1,L_SIZE),
				to_sfixed(-0.9922,1,L_SIZE),
				to_sfixed(-0.9922,1,L_SIZE),
				to_sfixed(-0.9922,1,L_SIZE),
				to_sfixed(-0.9922,1,L_SIZE),
				to_sfixed(-0.9922,1,L_SIZE),
				to_sfixed(-0.9921,1,L_SIZE),
				to_sfixed(-0.9921,1,L_SIZE),
				to_sfixed(-0.9921,1,L_SIZE),
				to_sfixed(-0.9921,1,L_SIZE),
				to_sfixed(-0.9921,1,L_SIZE),
				to_sfixed(-0.9921,1,L_SIZE),
				to_sfixed(-0.9921,1,L_SIZE),
				to_sfixed(-0.9921,1,L_SIZE),
				to_sfixed(-0.9921,1,L_SIZE),
				to_sfixed(-0.9921,1,L_SIZE),
				to_sfixed(-0.9921,1,L_SIZE),
				to_sfixed(-0.9921,1,L_SIZE),
				to_sfixed(-0.9921,1,L_SIZE),
				to_sfixed(-0.9921,1,L_SIZE),
				to_sfixed(-0.9921,1,L_SIZE),
				to_sfixed(-0.9921,1,L_SIZE),
				to_sfixed(-0.9921,1,L_SIZE),
				to_sfixed(-0.9921,1,L_SIZE),
				to_sfixed(-0.9920,1,L_SIZE),
				to_sfixed(-0.9920,1,L_SIZE),
				to_sfixed(-0.9920,1,L_SIZE),
				to_sfixed(-0.9920,1,L_SIZE),
				to_sfixed(-0.9920,1,L_SIZE),
				to_sfixed(-0.9920,1,L_SIZE),
				to_sfixed(-0.9920,1,L_SIZE),
				to_sfixed(-0.9920,1,L_SIZE),
				to_sfixed(-0.9920,1,L_SIZE),
				to_sfixed(-0.9920,1,L_SIZE),
				to_sfixed(-0.9920,1,L_SIZE),
				to_sfixed(-0.9920,1,L_SIZE),
				to_sfixed(-0.9920,1,L_SIZE),
				to_sfixed(-0.9920,1,L_SIZE),
				to_sfixed(-0.9920,1,L_SIZE),
				to_sfixed(-0.9920,1,L_SIZE),
				to_sfixed(-0.9920,1,L_SIZE),
				to_sfixed(-0.9919,1,L_SIZE),
				to_sfixed(-0.9919,1,L_SIZE),
				to_sfixed(-0.9919,1,L_SIZE),
				to_sfixed(-0.9919,1,L_SIZE),
				to_sfixed(-0.9919,1,L_SIZE),
				to_sfixed(-0.9919,1,L_SIZE),
				to_sfixed(-0.9919,1,L_SIZE),
				to_sfixed(-0.9919,1,L_SIZE),
				to_sfixed(-0.9919,1,L_SIZE),
				to_sfixed(-0.9919,1,L_SIZE),
				to_sfixed(-0.9919,1,L_SIZE),
				to_sfixed(-0.9919,1,L_SIZE),
				to_sfixed(-0.9919,1,L_SIZE),
				to_sfixed(-0.9919,1,L_SIZE),
				to_sfixed(-0.9919,1,L_SIZE),
				to_sfixed(-0.9919,1,L_SIZE),
				to_sfixed(-0.9919,1,L_SIZE),
				to_sfixed(-0.9918,1,L_SIZE),
				to_sfixed(-0.9918,1,L_SIZE),
				to_sfixed(-0.9918,1,L_SIZE),
				to_sfixed(-0.9918,1,L_SIZE),
				to_sfixed(-0.9918,1,L_SIZE),
				to_sfixed(-0.9918,1,L_SIZE),
				to_sfixed(-0.9918,1,L_SIZE),
				to_sfixed(-0.9918,1,L_SIZE),
				to_sfixed(-0.9918,1,L_SIZE),
				to_sfixed(-0.9918,1,L_SIZE),
				to_sfixed(-0.9918,1,L_SIZE),
				to_sfixed(-0.9918,1,L_SIZE),
				to_sfixed(-0.9918,1,L_SIZE),
				to_sfixed(-0.9918,1,L_SIZE),
				to_sfixed(-0.9918,1,L_SIZE),
				to_sfixed(-0.9918,1,L_SIZE),
				to_sfixed(-0.9918,1,L_SIZE),
				to_sfixed(-0.9917,1,L_SIZE),
				to_sfixed(-0.9917,1,L_SIZE),
				to_sfixed(-0.9917,1,L_SIZE),
				to_sfixed(-0.9917,1,L_SIZE),
				to_sfixed(-0.9917,1,L_SIZE),
				to_sfixed(-0.9917,1,L_SIZE),
				to_sfixed(-0.9917,1,L_SIZE),
				to_sfixed(-0.9917,1,L_SIZE),
				to_sfixed(-0.9917,1,L_SIZE),
				to_sfixed(-0.9917,1,L_SIZE),
				to_sfixed(-0.9917,1,L_SIZE),
				to_sfixed(-0.9917,1,L_SIZE),
				to_sfixed(-0.9917,1,L_SIZE),
				to_sfixed(-0.9917,1,L_SIZE),
				to_sfixed(-0.9917,1,L_SIZE),
				to_sfixed(-0.9917,1,L_SIZE),
				to_sfixed(-0.9916,1,L_SIZE),
				to_sfixed(-0.9916,1,L_SIZE),
				to_sfixed(-0.9916,1,L_SIZE),
				to_sfixed(-0.9916,1,L_SIZE),
				to_sfixed(-0.9916,1,L_SIZE),
				to_sfixed(-0.9916,1,L_SIZE),
				to_sfixed(-0.9916,1,L_SIZE),
				to_sfixed(-0.9916,1,L_SIZE),
				to_sfixed(-0.9916,1,L_SIZE),
				to_sfixed(-0.9916,1,L_SIZE),
				to_sfixed(-0.9916,1,L_SIZE),
				to_sfixed(-0.9916,1,L_SIZE),
				to_sfixed(-0.9916,1,L_SIZE),
				to_sfixed(-0.9916,1,L_SIZE),
				to_sfixed(-0.9916,1,L_SIZE),
				to_sfixed(-0.9916,1,L_SIZE),
				to_sfixed(-0.9915,1,L_SIZE),
				to_sfixed(-0.9915,1,L_SIZE),
				to_sfixed(-0.9915,1,L_SIZE),
				to_sfixed(-0.9915,1,L_SIZE),
				to_sfixed(-0.9915,1,L_SIZE),
				to_sfixed(-0.9915,1,L_SIZE),
				to_sfixed(-0.9915,1,L_SIZE),
				to_sfixed(-0.9915,1,L_SIZE),
				to_sfixed(-0.9915,1,L_SIZE),
				to_sfixed(-0.9915,1,L_SIZE),
				to_sfixed(-0.9915,1,L_SIZE),
				to_sfixed(-0.9915,1,L_SIZE),
				to_sfixed(-0.9915,1,L_SIZE),
				to_sfixed(-0.9915,1,L_SIZE),
				to_sfixed(-0.9915,1,L_SIZE),
				to_sfixed(-0.9915,1,L_SIZE),
				to_sfixed(-0.9914,1,L_SIZE),
				to_sfixed(-0.9914,1,L_SIZE),
				to_sfixed(-0.9914,1,L_SIZE),
				to_sfixed(-0.9914,1,L_SIZE),
				to_sfixed(-0.9914,1,L_SIZE),
				to_sfixed(-0.9914,1,L_SIZE),
				to_sfixed(-0.9914,1,L_SIZE),
				to_sfixed(-0.9914,1,L_SIZE),
				to_sfixed(-0.9914,1,L_SIZE),
				to_sfixed(-0.9914,1,L_SIZE),
				to_sfixed(-0.9914,1,L_SIZE),
				to_sfixed(-0.9914,1,L_SIZE),
				to_sfixed(-0.9914,1,L_SIZE),
				to_sfixed(-0.9914,1,L_SIZE),
				to_sfixed(-0.9914,1,L_SIZE),
				to_sfixed(-0.9914,1,L_SIZE),
				to_sfixed(-0.9913,1,L_SIZE),
				to_sfixed(-0.9913,1,L_SIZE),
				to_sfixed(-0.9913,1,L_SIZE),
				to_sfixed(-0.9913,1,L_SIZE),
				to_sfixed(-0.9913,1,L_SIZE),
				to_sfixed(-0.9913,1,L_SIZE),
				to_sfixed(-0.9913,1,L_SIZE),
				to_sfixed(-0.9913,1,L_SIZE),
				to_sfixed(-0.9913,1,L_SIZE),
				to_sfixed(-0.9913,1,L_SIZE),
				to_sfixed(-0.9913,1,L_SIZE),
				to_sfixed(-0.9913,1,L_SIZE),
				to_sfixed(-0.9913,1,L_SIZE),
				to_sfixed(-0.9913,1,L_SIZE),
				to_sfixed(-0.9913,1,L_SIZE),
				to_sfixed(-0.9913,1,L_SIZE),
				to_sfixed(-0.9912,1,L_SIZE),
				to_sfixed(-0.9912,1,L_SIZE),
				to_sfixed(-0.9912,1,L_SIZE),
				to_sfixed(-0.9912,1,L_SIZE),
				to_sfixed(-0.9912,1,L_SIZE),
				to_sfixed(-0.9912,1,L_SIZE),
				to_sfixed(-0.9912,1,L_SIZE),
				to_sfixed(-0.9912,1,L_SIZE),
				to_sfixed(-0.9912,1,L_SIZE),
				to_sfixed(-0.9912,1,L_SIZE),
				to_sfixed(-0.9912,1,L_SIZE),
				to_sfixed(-0.9912,1,L_SIZE),
				to_sfixed(-0.9912,1,L_SIZE),
				to_sfixed(-0.9912,1,L_SIZE),
				to_sfixed(-0.9912,1,L_SIZE),
				to_sfixed(-0.9912,1,L_SIZE),
				to_sfixed(-0.9911,1,L_SIZE),
				to_sfixed(-0.9911,1,L_SIZE),
				to_sfixed(-0.9911,1,L_SIZE),
				to_sfixed(-0.9911,1,L_SIZE),
				to_sfixed(-0.9911,1,L_SIZE),
				to_sfixed(-0.9911,1,L_SIZE),
				to_sfixed(-0.9911,1,L_SIZE),
				to_sfixed(-0.9911,1,L_SIZE),
				to_sfixed(-0.9911,1,L_SIZE),
				to_sfixed(-0.9911,1,L_SIZE),
				to_sfixed(-0.9911,1,L_SIZE),
				to_sfixed(-0.9911,1,L_SIZE),
				to_sfixed(-0.9911,1,L_SIZE),
				to_sfixed(-0.9911,1,L_SIZE),
				to_sfixed(-0.9911,1,L_SIZE),
				to_sfixed(-0.9910,1,L_SIZE),
				to_sfixed(-0.9910,1,L_SIZE),
				to_sfixed(-0.9910,1,L_SIZE),
				to_sfixed(-0.9910,1,L_SIZE),
				to_sfixed(-0.9910,1,L_SIZE),
				to_sfixed(-0.9910,1,L_SIZE),
				to_sfixed(-0.9910,1,L_SIZE),
				to_sfixed(-0.9910,1,L_SIZE),
				to_sfixed(-0.9910,1,L_SIZE),
				to_sfixed(-0.9910,1,L_SIZE),
				to_sfixed(-0.9910,1,L_SIZE),
				to_sfixed(-0.9910,1,L_SIZE),
				to_sfixed(-0.9910,1,L_SIZE),
				to_sfixed(-0.9910,1,L_SIZE),
				to_sfixed(-0.9910,1,L_SIZE),
				to_sfixed(-0.9909,1,L_SIZE),
				to_sfixed(-0.9909,1,L_SIZE),
				to_sfixed(-0.9909,1,L_SIZE),
				to_sfixed(-0.9909,1,L_SIZE),
				to_sfixed(-0.9909,1,L_SIZE),
				to_sfixed(-0.9909,1,L_SIZE),
				to_sfixed(-0.9909,1,L_SIZE),
				to_sfixed(-0.9909,1,L_SIZE),
				to_sfixed(-0.9909,1,L_SIZE),
				to_sfixed(-0.9909,1,L_SIZE),
				to_sfixed(-0.9909,1,L_SIZE),
				to_sfixed(-0.9909,1,L_SIZE),
				to_sfixed(-0.9909,1,L_SIZE),
				to_sfixed(-0.9909,1,L_SIZE),
				to_sfixed(-0.9909,1,L_SIZE),
				to_sfixed(-0.9909,1,L_SIZE),
				to_sfixed(-0.9908,1,L_SIZE),
				to_sfixed(-0.9908,1,L_SIZE),
				to_sfixed(-0.9908,1,L_SIZE),
				to_sfixed(-0.9908,1,L_SIZE),
				to_sfixed(-0.9908,1,L_SIZE),
				to_sfixed(-0.9908,1,L_SIZE),
				to_sfixed(-0.9908,1,L_SIZE),
				to_sfixed(-0.9908,1,L_SIZE),
				to_sfixed(-0.9908,1,L_SIZE),
				to_sfixed(-0.9908,1,L_SIZE),
				to_sfixed(-0.9908,1,L_SIZE),
				to_sfixed(-0.9908,1,L_SIZE),
				to_sfixed(-0.9908,1,L_SIZE),
				to_sfixed(-0.9908,1,L_SIZE),
				to_sfixed(-0.9907,1,L_SIZE),
				to_sfixed(-0.9907,1,L_SIZE),
				to_sfixed(-0.9907,1,L_SIZE),
				to_sfixed(-0.9907,1,L_SIZE),
				to_sfixed(-0.9907,1,L_SIZE),
				to_sfixed(-0.9907,1,L_SIZE),
				to_sfixed(-0.9907,1,L_SIZE),
				to_sfixed(-0.9907,1,L_SIZE),
				to_sfixed(-0.9907,1,L_SIZE),
				to_sfixed(-0.9907,1,L_SIZE),
				to_sfixed(-0.9907,1,L_SIZE),
				to_sfixed(-0.9907,1,L_SIZE),
				to_sfixed(-0.9907,1,L_SIZE),
				to_sfixed(-0.9907,1,L_SIZE),
				to_sfixed(-0.9907,1,L_SIZE),
				to_sfixed(-0.9906,1,L_SIZE),
				to_sfixed(-0.9906,1,L_SIZE),
				to_sfixed(-0.9906,1,L_SIZE),
				to_sfixed(-0.9906,1,L_SIZE),
				to_sfixed(-0.9906,1,L_SIZE),
				to_sfixed(-0.9906,1,L_SIZE),
				to_sfixed(-0.9906,1,L_SIZE),
				to_sfixed(-0.9906,1,L_SIZE),
				to_sfixed(-0.9906,1,L_SIZE),
				to_sfixed(-0.9906,1,L_SIZE),
				to_sfixed(-0.9906,1,L_SIZE),
				to_sfixed(-0.9906,1,L_SIZE),
				to_sfixed(-0.9906,1,L_SIZE),
				to_sfixed(-0.9906,1,L_SIZE),
				to_sfixed(-0.9906,1,L_SIZE),
				to_sfixed(-0.9905,1,L_SIZE),
				to_sfixed(-0.9905,1,L_SIZE),
				to_sfixed(-0.9905,1,L_SIZE),
				to_sfixed(-0.9905,1,L_SIZE),
				to_sfixed(-0.9905,1,L_SIZE),
				to_sfixed(-0.9905,1,L_SIZE),
				to_sfixed(-0.9905,1,L_SIZE),
				to_sfixed(-0.9905,1,L_SIZE),
				to_sfixed(-0.9905,1,L_SIZE),
				to_sfixed(-0.9905,1,L_SIZE),
				to_sfixed(-0.9905,1,L_SIZE),
				to_sfixed(-0.9905,1,L_SIZE),
				to_sfixed(-0.9905,1,L_SIZE),
				to_sfixed(-0.9905,1,L_SIZE),
				to_sfixed(-0.9904,1,L_SIZE),
				to_sfixed(-0.9904,1,L_SIZE),
				to_sfixed(-0.9904,1,L_SIZE),
				to_sfixed(-0.9904,1,L_SIZE),
				to_sfixed(-0.9904,1,L_SIZE),
				to_sfixed(-0.9904,1,L_SIZE),
				to_sfixed(-0.9904,1,L_SIZE),
				to_sfixed(-0.9904,1,L_SIZE),
				to_sfixed(-0.9904,1,L_SIZE),
				to_sfixed(-0.9904,1,L_SIZE),
				to_sfixed(-0.9904,1,L_SIZE),
				to_sfixed(-0.9904,1,L_SIZE),
				to_sfixed(-0.9904,1,L_SIZE),
				to_sfixed(-0.9904,1,L_SIZE),
				to_sfixed(-0.9903,1,L_SIZE),
				to_sfixed(-0.9903,1,L_SIZE),
				to_sfixed(-0.9903,1,L_SIZE),
				to_sfixed(-0.9903,1,L_SIZE),
				to_sfixed(-0.9903,1,L_SIZE),
				to_sfixed(-0.9903,1,L_SIZE),
				to_sfixed(-0.9903,1,L_SIZE),
				to_sfixed(-0.9903,1,L_SIZE),
				to_sfixed(-0.9903,1,L_SIZE),
				to_sfixed(-0.9903,1,L_SIZE),
				to_sfixed(-0.9903,1,L_SIZE),
				to_sfixed(-0.9903,1,L_SIZE),
				to_sfixed(-0.9903,1,L_SIZE),
				to_sfixed(-0.9903,1,L_SIZE),
				to_sfixed(-0.9903,1,L_SIZE),
				to_sfixed(-0.9902,1,L_SIZE),
				to_sfixed(-0.9902,1,L_SIZE),
				to_sfixed(-0.9902,1,L_SIZE),
				to_sfixed(-0.9902,1,L_SIZE),
				to_sfixed(-0.9902,1,L_SIZE),
				to_sfixed(-0.9902,1,L_SIZE),
				to_sfixed(-0.9902,1,L_SIZE),
				to_sfixed(-0.9902,1,L_SIZE),
				to_sfixed(-0.9902,1,L_SIZE),
				to_sfixed(-0.9902,1,L_SIZE),
				to_sfixed(-0.9902,1,L_SIZE),
				to_sfixed(-0.9902,1,L_SIZE),
				to_sfixed(-0.9902,1,L_SIZE),
				to_sfixed(-0.9902,1,L_SIZE),
				to_sfixed(-0.9901,1,L_SIZE),
				to_sfixed(-0.9901,1,L_SIZE),
				to_sfixed(-0.9901,1,L_SIZE),
				to_sfixed(-0.9901,1,L_SIZE),
				to_sfixed(-0.9901,1,L_SIZE),
				to_sfixed(-0.9901,1,L_SIZE),
				to_sfixed(-0.9901,1,L_SIZE),
				to_sfixed(-0.9901,1,L_SIZE),
				to_sfixed(-0.9901,1,L_SIZE),
				to_sfixed(-0.9901,1,L_SIZE),
				to_sfixed(-0.9901,1,L_SIZE),
				to_sfixed(-0.9901,1,L_SIZE),
				to_sfixed(-0.9901,1,L_SIZE),
				to_sfixed(-0.9900,1,L_SIZE),
				to_sfixed(-0.9900,1,L_SIZE),
				to_sfixed(-0.9900,1,L_SIZE),
				to_sfixed(-0.9900,1,L_SIZE),
				to_sfixed(-0.9900,1,L_SIZE),
				to_sfixed(-0.9900,1,L_SIZE),
				to_sfixed(-0.9900,1,L_SIZE),
				to_sfixed(-0.9900,1,L_SIZE),
				to_sfixed(-0.9900,1,L_SIZE),
				to_sfixed(-0.9900,1,L_SIZE),
				to_sfixed(-0.9900,1,L_SIZE),
				to_sfixed(-0.9900,1,L_SIZE),
				to_sfixed(-0.9900,1,L_SIZE),
				to_sfixed(-0.9900,1,L_SIZE),
				to_sfixed(-0.9899,1,L_SIZE),
				to_sfixed(-0.9899,1,L_SIZE),
				to_sfixed(-0.9899,1,L_SIZE),
				to_sfixed(-0.9899,1,L_SIZE),
				to_sfixed(-0.9899,1,L_SIZE),
				to_sfixed(-0.9899,1,L_SIZE),
				to_sfixed(-0.9899,1,L_SIZE),
				to_sfixed(-0.9899,1,L_SIZE),
				to_sfixed(-0.9899,1,L_SIZE),
				to_sfixed(-0.9899,1,L_SIZE),
				to_sfixed(-0.9899,1,L_SIZE),
				to_sfixed(-0.9899,1,L_SIZE),
				to_sfixed(-0.9899,1,L_SIZE),
				to_sfixed(-0.9899,1,L_SIZE),
				to_sfixed(-0.9898,1,L_SIZE),
				to_sfixed(-0.9898,1,L_SIZE),
				to_sfixed(-0.9898,1,L_SIZE),
				to_sfixed(-0.9898,1,L_SIZE),
				to_sfixed(-0.9898,1,L_SIZE),
				to_sfixed(-0.9898,1,L_SIZE),
				to_sfixed(-0.9898,1,L_SIZE),
				to_sfixed(-0.9898,1,L_SIZE),
				to_sfixed(-0.9898,1,L_SIZE),
				to_sfixed(-0.9898,1,L_SIZE),
				to_sfixed(-0.9898,1,L_SIZE),
				to_sfixed(-0.9898,1,L_SIZE),
				to_sfixed(-0.9898,1,L_SIZE),
				to_sfixed(-0.9897,1,L_SIZE),
				to_sfixed(-0.9897,1,L_SIZE),
				to_sfixed(-0.9897,1,L_SIZE),
				to_sfixed(-0.9897,1,L_SIZE),
				to_sfixed(-0.9897,1,L_SIZE),
				to_sfixed(-0.9897,1,L_SIZE),
				to_sfixed(-0.9897,1,L_SIZE),
				to_sfixed(-0.9897,1,L_SIZE),
				to_sfixed(-0.9897,1,L_SIZE),
				to_sfixed(-0.9897,1,L_SIZE),
				to_sfixed(-0.9897,1,L_SIZE),
				to_sfixed(-0.9897,1,L_SIZE),
				to_sfixed(-0.9897,1,L_SIZE),
				to_sfixed(-0.9897,1,L_SIZE),
				to_sfixed(-0.9896,1,L_SIZE),
				to_sfixed(-0.9896,1,L_SIZE),
				to_sfixed(-0.9896,1,L_SIZE),
				to_sfixed(-0.9896,1,L_SIZE),
				to_sfixed(-0.9896,1,L_SIZE),
				to_sfixed(-0.9896,1,L_SIZE),
				to_sfixed(-0.9896,1,L_SIZE),
				to_sfixed(-0.9896,1,L_SIZE),
				to_sfixed(-0.9896,1,L_SIZE),
				to_sfixed(-0.9896,1,L_SIZE),
				to_sfixed(-0.9896,1,L_SIZE),
				to_sfixed(-0.9896,1,L_SIZE),
				to_sfixed(-0.9896,1,L_SIZE),
				to_sfixed(-0.9895,1,L_SIZE),
				to_sfixed(-0.9895,1,L_SIZE),
				to_sfixed(-0.9895,1,L_SIZE),
				to_sfixed(-0.9895,1,L_SIZE),
				to_sfixed(-0.9895,1,L_SIZE),
				to_sfixed(-0.9895,1,L_SIZE),
				to_sfixed(-0.9895,1,L_SIZE),
				to_sfixed(-0.9895,1,L_SIZE),
				to_sfixed(-0.9895,1,L_SIZE),
				to_sfixed(-0.9895,1,L_SIZE),
				to_sfixed(-0.9895,1,L_SIZE),
				to_sfixed(-0.9895,1,L_SIZE),
				to_sfixed(-0.9895,1,L_SIZE),
				to_sfixed(-0.9894,1,L_SIZE),
				to_sfixed(-0.9894,1,L_SIZE),
				to_sfixed(-0.9894,1,L_SIZE),
				to_sfixed(-0.9894,1,L_SIZE),
				to_sfixed(-0.9894,1,L_SIZE),
				to_sfixed(-0.9894,1,L_SIZE),
				to_sfixed(-0.9894,1,L_SIZE),
				to_sfixed(-0.9894,1,L_SIZE),
				to_sfixed(-0.9894,1,L_SIZE),
				to_sfixed(-0.9894,1,L_SIZE),
				to_sfixed(-0.9894,1,L_SIZE),
				to_sfixed(-0.9894,1,L_SIZE),
				to_sfixed(-0.9894,1,L_SIZE),
				to_sfixed(-0.9893,1,L_SIZE),
				to_sfixed(-0.9893,1,L_SIZE),
				to_sfixed(-0.9893,1,L_SIZE),
				to_sfixed(-0.9893,1,L_SIZE),
				to_sfixed(-0.9893,1,L_SIZE),
				to_sfixed(-0.9893,1,L_SIZE),
				to_sfixed(-0.9893,1,L_SIZE),
				to_sfixed(-0.9893,1,L_SIZE),
				to_sfixed(-0.9893,1,L_SIZE),
				to_sfixed(-0.9893,1,L_SIZE),
				to_sfixed(-0.9893,1,L_SIZE),
				to_sfixed(-0.9893,1,L_SIZE),
				to_sfixed(-0.9893,1,L_SIZE),
				to_sfixed(-0.9892,1,L_SIZE),
				to_sfixed(-0.9892,1,L_SIZE),
				to_sfixed(-0.9892,1,L_SIZE),
				to_sfixed(-0.9892,1,L_SIZE),
				to_sfixed(-0.9892,1,L_SIZE),
				to_sfixed(-0.9892,1,L_SIZE),
				to_sfixed(-0.9892,1,L_SIZE),
				to_sfixed(-0.9892,1,L_SIZE),
				to_sfixed(-0.9892,1,L_SIZE),
				to_sfixed(-0.9892,1,L_SIZE),
				to_sfixed(-0.9892,1,L_SIZE),
				to_sfixed(-0.9892,1,L_SIZE),
				to_sfixed(-0.9891,1,L_SIZE),
				to_sfixed(-0.9891,1,L_SIZE),
				to_sfixed(-0.9891,1,L_SIZE),
				to_sfixed(-0.9891,1,L_SIZE),
				to_sfixed(-0.9891,1,L_SIZE),
				to_sfixed(-0.9891,1,L_SIZE),
				to_sfixed(-0.9891,1,L_SIZE),
				to_sfixed(-0.9891,1,L_SIZE),
				to_sfixed(-0.9891,1,L_SIZE),
				to_sfixed(-0.9891,1,L_SIZE),
				to_sfixed(-0.9891,1,L_SIZE),
				to_sfixed(-0.9891,1,L_SIZE),
				to_sfixed(-0.9891,1,L_SIZE),
				to_sfixed(-0.9890,1,L_SIZE),
				to_sfixed(-0.9890,1,L_SIZE),
				to_sfixed(-0.9890,1,L_SIZE),
				to_sfixed(-0.9890,1,L_SIZE),
				to_sfixed(-0.9890,1,L_SIZE),
				to_sfixed(-0.9890,1,L_SIZE),
				to_sfixed(-0.9890,1,L_SIZE),
				to_sfixed(-0.9890,1,L_SIZE),
				to_sfixed(-0.9890,1,L_SIZE),
				to_sfixed(-0.9890,1,L_SIZE),
				to_sfixed(-0.9890,1,L_SIZE),
				to_sfixed(-0.9890,1,L_SIZE),
				to_sfixed(-0.9889,1,L_SIZE),
				to_sfixed(-0.9889,1,L_SIZE),
				to_sfixed(-0.9889,1,L_SIZE),
				to_sfixed(-0.9889,1,L_SIZE),
				to_sfixed(-0.9889,1,L_SIZE),
				to_sfixed(-0.9889,1,L_SIZE),
				to_sfixed(-0.9889,1,L_SIZE),
				to_sfixed(-0.9889,1,L_SIZE),
				to_sfixed(-0.9889,1,L_SIZE),
				to_sfixed(-0.9889,1,L_SIZE),
				to_sfixed(-0.9889,1,L_SIZE),
				to_sfixed(-0.9889,1,L_SIZE),
				to_sfixed(-0.9889,1,L_SIZE),
				to_sfixed(-0.9888,1,L_SIZE),
				to_sfixed(-0.9888,1,L_SIZE),
				to_sfixed(-0.9888,1,L_SIZE),
				to_sfixed(-0.9888,1,L_SIZE),
				to_sfixed(-0.9888,1,L_SIZE),
				to_sfixed(-0.9888,1,L_SIZE),
				to_sfixed(-0.9888,1,L_SIZE),
				to_sfixed(-0.9888,1,L_SIZE),
				to_sfixed(-0.9888,1,L_SIZE),
				to_sfixed(-0.9888,1,L_SIZE),
				to_sfixed(-0.9888,1,L_SIZE),
				to_sfixed(-0.9888,1,L_SIZE),
				to_sfixed(-0.9887,1,L_SIZE),
				to_sfixed(-0.9887,1,L_SIZE),
				to_sfixed(-0.9887,1,L_SIZE),
				to_sfixed(-0.9887,1,L_SIZE),
				to_sfixed(-0.9887,1,L_SIZE),
				to_sfixed(-0.9887,1,L_SIZE),
				to_sfixed(-0.9887,1,L_SIZE),
				to_sfixed(-0.9887,1,L_SIZE),
				to_sfixed(-0.9887,1,L_SIZE),
				to_sfixed(-0.9887,1,L_SIZE),
				to_sfixed(-0.9887,1,L_SIZE),
				to_sfixed(-0.9887,1,L_SIZE),
				to_sfixed(-0.9886,1,L_SIZE),
				to_sfixed(-0.9886,1,L_SIZE),
				to_sfixed(-0.9886,1,L_SIZE),
				to_sfixed(-0.9886,1,L_SIZE),
				to_sfixed(-0.9886,1,L_SIZE),
				to_sfixed(-0.9886,1,L_SIZE),
				to_sfixed(-0.9886,1,L_SIZE),
				to_sfixed(-0.9886,1,L_SIZE),
				to_sfixed(-0.9886,1,L_SIZE),
				to_sfixed(-0.9886,1,L_SIZE),
				to_sfixed(-0.9886,1,L_SIZE),
				to_sfixed(-0.9886,1,L_SIZE),
				to_sfixed(-0.9885,1,L_SIZE),
				to_sfixed(-0.9885,1,L_SIZE),
				to_sfixed(-0.9885,1,L_SIZE),
				to_sfixed(-0.9885,1,L_SIZE),
				to_sfixed(-0.9885,1,L_SIZE),
				to_sfixed(-0.9885,1,L_SIZE),
				to_sfixed(-0.9885,1,L_SIZE),
				to_sfixed(-0.9885,1,L_SIZE),
				to_sfixed(-0.9885,1,L_SIZE),
				to_sfixed(-0.9885,1,L_SIZE),
				to_sfixed(-0.9885,1,L_SIZE),
				to_sfixed(-0.9885,1,L_SIZE),
				to_sfixed(-0.9884,1,L_SIZE),
				to_sfixed(-0.9884,1,L_SIZE),
				to_sfixed(-0.9884,1,L_SIZE),
				to_sfixed(-0.9884,1,L_SIZE),
				to_sfixed(-0.9884,1,L_SIZE),
				to_sfixed(-0.9884,1,L_SIZE),
				to_sfixed(-0.9884,1,L_SIZE),
				to_sfixed(-0.9884,1,L_SIZE),
				to_sfixed(-0.9884,1,L_SIZE),
				to_sfixed(-0.9884,1,L_SIZE),
				to_sfixed(-0.9884,1,L_SIZE),
				to_sfixed(-0.9884,1,L_SIZE),
				to_sfixed(-0.9883,1,L_SIZE),
				to_sfixed(-0.9883,1,L_SIZE),
				to_sfixed(-0.9883,1,L_SIZE),
				to_sfixed(-0.9883,1,L_SIZE),
				to_sfixed(-0.9883,1,L_SIZE),
				to_sfixed(-0.9883,1,L_SIZE),
				to_sfixed(-0.9883,1,L_SIZE),
				to_sfixed(-0.9883,1,L_SIZE),
				to_sfixed(-0.9883,1,L_SIZE),
				to_sfixed(-0.9883,1,L_SIZE),
				to_sfixed(-0.9883,1,L_SIZE),
				to_sfixed(-0.9883,1,L_SIZE),
				to_sfixed(-0.9882,1,L_SIZE),
				to_sfixed(-0.9882,1,L_SIZE),
				to_sfixed(-0.9882,1,L_SIZE),
				to_sfixed(-0.9882,1,L_SIZE),
				to_sfixed(-0.9882,1,L_SIZE),
				to_sfixed(-0.9882,1,L_SIZE),
				to_sfixed(-0.9882,1,L_SIZE),
				to_sfixed(-0.9882,1,L_SIZE),
				to_sfixed(-0.9882,1,L_SIZE),
				to_sfixed(-0.9882,1,L_SIZE),
				to_sfixed(-0.9882,1,L_SIZE),
				to_sfixed(-0.9881,1,L_SIZE),
				to_sfixed(-0.9881,1,L_SIZE),
				to_sfixed(-0.9881,1,L_SIZE),
				to_sfixed(-0.9881,1,L_SIZE),
				to_sfixed(-0.9881,1,L_SIZE),
				to_sfixed(-0.9881,1,L_SIZE),
				to_sfixed(-0.9881,1,L_SIZE),
				to_sfixed(-0.9881,1,L_SIZE),
				to_sfixed(-0.9881,1,L_SIZE),
				to_sfixed(-0.9881,1,L_SIZE),
				to_sfixed(-0.9881,1,L_SIZE),
				to_sfixed(-0.9881,1,L_SIZE),
				to_sfixed(-0.9880,1,L_SIZE),
				to_sfixed(-0.9880,1,L_SIZE),
				to_sfixed(-0.9880,1,L_SIZE),
				to_sfixed(-0.9880,1,L_SIZE),
				to_sfixed(-0.9880,1,L_SIZE),
				to_sfixed(-0.9880,1,L_SIZE),
				to_sfixed(-0.9880,1,L_SIZE),
				to_sfixed(-0.9880,1,L_SIZE),
				to_sfixed(-0.9880,1,L_SIZE),
				to_sfixed(-0.9880,1,L_SIZE),
				to_sfixed(-0.9880,1,L_SIZE),
				to_sfixed(-0.9879,1,L_SIZE),
				to_sfixed(-0.9879,1,L_SIZE),
				to_sfixed(-0.9879,1,L_SIZE),
				to_sfixed(-0.9879,1,L_SIZE),
				to_sfixed(-0.9879,1,L_SIZE),
				to_sfixed(-0.9879,1,L_SIZE),
				to_sfixed(-0.9879,1,L_SIZE),
				to_sfixed(-0.9879,1,L_SIZE),
				to_sfixed(-0.9879,1,L_SIZE),
				to_sfixed(-0.9879,1,L_SIZE),
				to_sfixed(-0.9879,1,L_SIZE),
				to_sfixed(-0.9879,1,L_SIZE),
				to_sfixed(-0.9878,1,L_SIZE),
				to_sfixed(-0.9878,1,L_SIZE),
				to_sfixed(-0.9878,1,L_SIZE),
				to_sfixed(-0.9878,1,L_SIZE),
				to_sfixed(-0.9878,1,L_SIZE),
				to_sfixed(-0.9878,1,L_SIZE),
				to_sfixed(-0.9878,1,L_SIZE),
				to_sfixed(-0.9878,1,L_SIZE),
				to_sfixed(-0.9878,1,L_SIZE),
				to_sfixed(-0.9878,1,L_SIZE),
				to_sfixed(-0.9878,1,L_SIZE),
				to_sfixed(-0.9877,1,L_SIZE),
				to_sfixed(-0.9877,1,L_SIZE),
				to_sfixed(-0.9877,1,L_SIZE),
				to_sfixed(-0.9877,1,L_SIZE),
				to_sfixed(-0.9877,1,L_SIZE),
				to_sfixed(-0.9877,1,L_SIZE),
				to_sfixed(-0.9877,1,L_SIZE),
				to_sfixed(-0.9877,1,L_SIZE),
				to_sfixed(-0.9877,1,L_SIZE),
				to_sfixed(-0.9877,1,L_SIZE),
				to_sfixed(-0.9877,1,L_SIZE),
				to_sfixed(-0.9876,1,L_SIZE),
				to_sfixed(-0.9876,1,L_SIZE),
				to_sfixed(-0.9876,1,L_SIZE),
				to_sfixed(-0.9876,1,L_SIZE),
				to_sfixed(-0.9876,1,L_SIZE),
				to_sfixed(-0.9876,1,L_SIZE),
				to_sfixed(-0.9876,1,L_SIZE),
				to_sfixed(-0.9876,1,L_SIZE),
				to_sfixed(-0.9876,1,L_SIZE),
				to_sfixed(-0.9876,1,L_SIZE),
				to_sfixed(-0.9876,1,L_SIZE),
				to_sfixed(-0.9875,1,L_SIZE),
				to_sfixed(-0.9875,1,L_SIZE),
				to_sfixed(-0.9875,1,L_SIZE),
				to_sfixed(-0.9875,1,L_SIZE),
				to_sfixed(-0.9875,1,L_SIZE),
				to_sfixed(-0.9875,1,L_SIZE),
				to_sfixed(-0.9875,1,L_SIZE),
				to_sfixed(-0.9875,1,L_SIZE),
				to_sfixed(-0.9875,1,L_SIZE),
				to_sfixed(-0.9875,1,L_SIZE),
				to_sfixed(-0.9875,1,L_SIZE),
				to_sfixed(-0.9874,1,L_SIZE),
				to_sfixed(-0.9874,1,L_SIZE),
				to_sfixed(-0.9874,1,L_SIZE),
				to_sfixed(-0.9874,1,L_SIZE),
				to_sfixed(-0.9874,1,L_SIZE),
				to_sfixed(-0.9874,1,L_SIZE),
				to_sfixed(-0.9874,1,L_SIZE),
				to_sfixed(-0.9874,1,L_SIZE),
				to_sfixed(-0.9874,1,L_SIZE),
				to_sfixed(-0.9874,1,L_SIZE),
				to_sfixed(-0.9874,1,L_SIZE),
				to_sfixed(-0.9873,1,L_SIZE),
				to_sfixed(-0.9873,1,L_SIZE),
				to_sfixed(-0.9873,1,L_SIZE),
				to_sfixed(-0.9873,1,L_SIZE),
				to_sfixed(-0.9873,1,L_SIZE),
				to_sfixed(-0.9873,1,L_SIZE),
				to_sfixed(-0.9873,1,L_SIZE),
				to_sfixed(-0.9873,1,L_SIZE),
				to_sfixed(-0.9873,1,L_SIZE),
				to_sfixed(-0.9873,1,L_SIZE),
				to_sfixed(-0.9873,1,L_SIZE),
				to_sfixed(-0.9872,1,L_SIZE),
				to_sfixed(-0.9872,1,L_SIZE),
				to_sfixed(-0.9872,1,L_SIZE),
				to_sfixed(-0.9872,1,L_SIZE),
				to_sfixed(-0.9872,1,L_SIZE),
				to_sfixed(-0.9872,1,L_SIZE),
				to_sfixed(-0.9872,1,L_SIZE),
				to_sfixed(-0.9872,1,L_SIZE),
				to_sfixed(-0.9872,1,L_SIZE),
				to_sfixed(-0.9872,1,L_SIZE),
				to_sfixed(-0.9872,1,L_SIZE),
				to_sfixed(-0.9871,1,L_SIZE),
				to_sfixed(-0.9871,1,L_SIZE),
				to_sfixed(-0.9871,1,L_SIZE),
				to_sfixed(-0.9871,1,L_SIZE),
				to_sfixed(-0.9871,1,L_SIZE),
				to_sfixed(-0.9871,1,L_SIZE),
				to_sfixed(-0.9871,1,L_SIZE),
				to_sfixed(-0.9871,1,L_SIZE),
				to_sfixed(-0.9871,1,L_SIZE),
				to_sfixed(-0.9871,1,L_SIZE),
				to_sfixed(-0.9870,1,L_SIZE),
				to_sfixed(-0.9870,1,L_SIZE),
				to_sfixed(-0.9870,1,L_SIZE),
				to_sfixed(-0.9870,1,L_SIZE),
				to_sfixed(-0.9870,1,L_SIZE),
				to_sfixed(-0.9870,1,L_SIZE),
				to_sfixed(-0.9870,1,L_SIZE),
				to_sfixed(-0.9870,1,L_SIZE),
				to_sfixed(-0.9870,1,L_SIZE),
				to_sfixed(-0.9870,1,L_SIZE),
				to_sfixed(-0.9870,1,L_SIZE),
				to_sfixed(-0.9869,1,L_SIZE),
				to_sfixed(-0.9869,1,L_SIZE),
				to_sfixed(-0.9869,1,L_SIZE),
				to_sfixed(-0.9869,1,L_SIZE),
				to_sfixed(-0.9869,1,L_SIZE),
				to_sfixed(-0.9869,1,L_SIZE),
				to_sfixed(-0.9869,1,L_SIZE),
				to_sfixed(-0.9869,1,L_SIZE),
				to_sfixed(-0.9869,1,L_SIZE),
				to_sfixed(-0.9869,1,L_SIZE),
				to_sfixed(-0.9868,1,L_SIZE),
				to_sfixed(-0.9868,1,L_SIZE),
				to_sfixed(-0.9868,1,L_SIZE),
				to_sfixed(-0.9868,1,L_SIZE),
				to_sfixed(-0.9868,1,L_SIZE),
				to_sfixed(-0.9868,1,L_SIZE),
				to_sfixed(-0.9868,1,L_SIZE),
				to_sfixed(-0.9868,1,L_SIZE),
				to_sfixed(-0.9868,1,L_SIZE),
				to_sfixed(-0.9868,1,L_SIZE),
				to_sfixed(-0.9868,1,L_SIZE),
				to_sfixed(-0.9867,1,L_SIZE),
				to_sfixed(-0.9867,1,L_SIZE),
				to_sfixed(-0.9867,1,L_SIZE),
				to_sfixed(-0.9867,1,L_SIZE),
				to_sfixed(-0.9867,1,L_SIZE),
				to_sfixed(-0.9867,1,L_SIZE),
				to_sfixed(-0.9867,1,L_SIZE),
				to_sfixed(-0.9867,1,L_SIZE),
				to_sfixed(-0.9867,1,L_SIZE),
				to_sfixed(-0.9867,1,L_SIZE),
				to_sfixed(-0.9866,1,L_SIZE),
				to_sfixed(-0.9866,1,L_SIZE),
				to_sfixed(-0.9866,1,L_SIZE),
				to_sfixed(-0.9866,1,L_SIZE),
				to_sfixed(-0.9866,1,L_SIZE),
				to_sfixed(-0.9866,1,L_SIZE),
				to_sfixed(-0.9866,1,L_SIZE),
				to_sfixed(-0.9866,1,L_SIZE),
				to_sfixed(-0.9866,1,L_SIZE),
				to_sfixed(-0.9866,1,L_SIZE),
				to_sfixed(-0.9865,1,L_SIZE),
				to_sfixed(-0.9865,1,L_SIZE),
				to_sfixed(-0.9865,1,L_SIZE),
				to_sfixed(-0.9865,1,L_SIZE),
				to_sfixed(-0.9865,1,L_SIZE),
				to_sfixed(-0.9865,1,L_SIZE),
				to_sfixed(-0.9865,1,L_SIZE),
				to_sfixed(-0.9865,1,L_SIZE),
				to_sfixed(-0.9865,1,L_SIZE),
				to_sfixed(-0.9865,1,L_SIZE),
				to_sfixed(-0.9865,1,L_SIZE),
				to_sfixed(-0.9864,1,L_SIZE),
				to_sfixed(-0.9864,1,L_SIZE),
				to_sfixed(-0.9864,1,L_SIZE),
				to_sfixed(-0.9864,1,L_SIZE),
				to_sfixed(-0.9864,1,L_SIZE),
				to_sfixed(-0.9864,1,L_SIZE),
				to_sfixed(-0.9864,1,L_SIZE),
				to_sfixed(-0.9864,1,L_SIZE),
				to_sfixed(-0.9864,1,L_SIZE),
				to_sfixed(-0.9864,1,L_SIZE),
				to_sfixed(-0.9863,1,L_SIZE),
				to_sfixed(-0.9863,1,L_SIZE),
				to_sfixed(-0.9863,1,L_SIZE),
				to_sfixed(-0.9863,1,L_SIZE),
				to_sfixed(-0.9863,1,L_SIZE),
				to_sfixed(-0.9863,1,L_SIZE),
				to_sfixed(-0.9863,1,L_SIZE),
				to_sfixed(-0.9863,1,L_SIZE),
				to_sfixed(-0.9863,1,L_SIZE),
				to_sfixed(-0.9863,1,L_SIZE),
				to_sfixed(-0.9862,1,L_SIZE),
				to_sfixed(-0.9862,1,L_SIZE),
				to_sfixed(-0.9862,1,L_SIZE),
				to_sfixed(-0.9862,1,L_SIZE),
				to_sfixed(-0.9862,1,L_SIZE),
				to_sfixed(-0.9862,1,L_SIZE),
				to_sfixed(-0.9862,1,L_SIZE),
				to_sfixed(-0.9862,1,L_SIZE),
				to_sfixed(-0.9862,1,L_SIZE),
				to_sfixed(-0.9862,1,L_SIZE),
				to_sfixed(-0.9861,1,L_SIZE),
				to_sfixed(-0.9861,1,L_SIZE),
				to_sfixed(-0.9861,1,L_SIZE),
				to_sfixed(-0.9861,1,L_SIZE),
				to_sfixed(-0.9861,1,L_SIZE),
				to_sfixed(-0.9861,1,L_SIZE),
				to_sfixed(-0.9861,1,L_SIZE),
				to_sfixed(-0.9861,1,L_SIZE),
				to_sfixed(-0.9861,1,L_SIZE),
				to_sfixed(-0.9861,1,L_SIZE),
				to_sfixed(-0.9860,1,L_SIZE),
				to_sfixed(-0.9860,1,L_SIZE),
				to_sfixed(-0.9860,1,L_SIZE),
				to_sfixed(-0.9860,1,L_SIZE),
				to_sfixed(-0.9860,1,L_SIZE),
				to_sfixed(-0.9860,1,L_SIZE),
				to_sfixed(-0.9860,1,L_SIZE),
				to_sfixed(-0.9860,1,L_SIZE),
				to_sfixed(-0.9860,1,L_SIZE),
				to_sfixed(-0.9859,1,L_SIZE),
				to_sfixed(-0.9859,1,L_SIZE),
				to_sfixed(-0.9859,1,L_SIZE),
				to_sfixed(-0.9859,1,L_SIZE),
				to_sfixed(-0.9859,1,L_SIZE),
				to_sfixed(-0.9859,1,L_SIZE),
				to_sfixed(-0.9859,1,L_SIZE),
				to_sfixed(-0.9859,1,L_SIZE),
				to_sfixed(-0.9859,1,L_SIZE),
				to_sfixed(-0.9859,1,L_SIZE),
				to_sfixed(-0.9858,1,L_SIZE),
				to_sfixed(-0.9858,1,L_SIZE),
				to_sfixed(-0.9858,1,L_SIZE),
				to_sfixed(-0.9858,1,L_SIZE),
				to_sfixed(-0.9858,1,L_SIZE),
				to_sfixed(-0.9858,1,L_SIZE),
				to_sfixed(-0.9858,1,L_SIZE),
				to_sfixed(-0.9858,1,L_SIZE),
				to_sfixed(-0.9858,1,L_SIZE),
				to_sfixed(-0.9858,1,L_SIZE),
				to_sfixed(-0.9857,1,L_SIZE),
				to_sfixed(-0.9857,1,L_SIZE),
				to_sfixed(-0.9857,1,L_SIZE),
				to_sfixed(-0.9857,1,L_SIZE),
				to_sfixed(-0.9857,1,L_SIZE),
				to_sfixed(-0.9857,1,L_SIZE),
				to_sfixed(-0.9857,1,L_SIZE),
				to_sfixed(-0.9857,1,L_SIZE),
				to_sfixed(-0.9857,1,L_SIZE),
				to_sfixed(-0.9856,1,L_SIZE),
				to_sfixed(-0.9856,1,L_SIZE),
				to_sfixed(-0.9856,1,L_SIZE),
				to_sfixed(-0.9856,1,L_SIZE),
				to_sfixed(-0.9856,1,L_SIZE),
				to_sfixed(-0.9856,1,L_SIZE),
				to_sfixed(-0.9856,1,L_SIZE),
				to_sfixed(-0.9856,1,L_SIZE),
				to_sfixed(-0.9856,1,L_SIZE),
				to_sfixed(-0.9856,1,L_SIZE),
				to_sfixed(-0.9855,1,L_SIZE),
				to_sfixed(-0.9855,1,L_SIZE),
				to_sfixed(-0.9855,1,L_SIZE),
				to_sfixed(-0.9855,1,L_SIZE),
				to_sfixed(-0.9855,1,L_SIZE),
				to_sfixed(-0.9855,1,L_SIZE),
				to_sfixed(-0.9855,1,L_SIZE),
				to_sfixed(-0.9855,1,L_SIZE),
				to_sfixed(-0.9855,1,L_SIZE),
				to_sfixed(-0.9855,1,L_SIZE),
				to_sfixed(-0.9854,1,L_SIZE),
				to_sfixed(-0.9854,1,L_SIZE),
				to_sfixed(-0.9854,1,L_SIZE),
				to_sfixed(-0.9854,1,L_SIZE),
				to_sfixed(-0.9854,1,L_SIZE),
				to_sfixed(-0.9854,1,L_SIZE),
				to_sfixed(-0.9854,1,L_SIZE),
				to_sfixed(-0.9854,1,L_SIZE),
				to_sfixed(-0.9854,1,L_SIZE),
				to_sfixed(-0.9853,1,L_SIZE),
				to_sfixed(-0.9853,1,L_SIZE),
				to_sfixed(-0.9853,1,L_SIZE),
				to_sfixed(-0.9853,1,L_SIZE),
				to_sfixed(-0.9853,1,L_SIZE),
				to_sfixed(-0.9853,1,L_SIZE),
				to_sfixed(-0.9853,1,L_SIZE),
				to_sfixed(-0.9853,1,L_SIZE),
				to_sfixed(-0.9853,1,L_SIZE),
				to_sfixed(-0.9852,1,L_SIZE),
				to_sfixed(-0.9852,1,L_SIZE),
				to_sfixed(-0.9852,1,L_SIZE),
				to_sfixed(-0.9852,1,L_SIZE),
				to_sfixed(-0.9852,1,L_SIZE),
				to_sfixed(-0.9852,1,L_SIZE),
				to_sfixed(-0.9852,1,L_SIZE),
				to_sfixed(-0.9852,1,L_SIZE),
				to_sfixed(-0.9852,1,L_SIZE),
				to_sfixed(-0.9852,1,L_SIZE),
				to_sfixed(-0.9851,1,L_SIZE),
				to_sfixed(-0.9851,1,L_SIZE),
				to_sfixed(-0.9851,1,L_SIZE),
				to_sfixed(-0.9851,1,L_SIZE),
				to_sfixed(-0.9851,1,L_SIZE),
				to_sfixed(-0.9851,1,L_SIZE),
				to_sfixed(-0.9851,1,L_SIZE),
				to_sfixed(-0.9851,1,L_SIZE),
				to_sfixed(-0.9851,1,L_SIZE),
				to_sfixed(-0.9850,1,L_SIZE),
				to_sfixed(-0.9850,1,L_SIZE),
				to_sfixed(-0.9850,1,L_SIZE),
				to_sfixed(-0.9850,1,L_SIZE),
				to_sfixed(-0.9850,1,L_SIZE),
				to_sfixed(-0.9850,1,L_SIZE),
				to_sfixed(-0.9850,1,L_SIZE),
				to_sfixed(-0.9850,1,L_SIZE),
				to_sfixed(-0.9850,1,L_SIZE),
				to_sfixed(-0.9849,1,L_SIZE),
				to_sfixed(-0.9849,1,L_SIZE),
				to_sfixed(-0.9849,1,L_SIZE),
				to_sfixed(-0.9849,1,L_SIZE),
				to_sfixed(-0.9849,1,L_SIZE),
				to_sfixed(-0.9849,1,L_SIZE),
				to_sfixed(-0.9849,1,L_SIZE),
				to_sfixed(-0.9849,1,L_SIZE),
				to_sfixed(-0.9849,1,L_SIZE),
				to_sfixed(-0.9848,1,L_SIZE),
				to_sfixed(-0.9848,1,L_SIZE),
				to_sfixed(-0.9848,1,L_SIZE),
				to_sfixed(-0.9848,1,L_SIZE),
				to_sfixed(-0.9848,1,L_SIZE),
				to_sfixed(-0.9848,1,L_SIZE),
				to_sfixed(-0.9848,1,L_SIZE),
				to_sfixed(-0.9848,1,L_SIZE),
				to_sfixed(-0.9848,1,L_SIZE),
				to_sfixed(-0.9847,1,L_SIZE),
				to_sfixed(-0.9847,1,L_SIZE),
				to_sfixed(-0.9847,1,L_SIZE),
				to_sfixed(-0.9847,1,L_SIZE),
				to_sfixed(-0.9847,1,L_SIZE),
				to_sfixed(-0.9847,1,L_SIZE),
				to_sfixed(-0.9847,1,L_SIZE),
				to_sfixed(-0.9847,1,L_SIZE),
				to_sfixed(-0.9847,1,L_SIZE),
				to_sfixed(-0.9846,1,L_SIZE),
				to_sfixed(-0.9846,1,L_SIZE),
				to_sfixed(-0.9846,1,L_SIZE),
				to_sfixed(-0.9846,1,L_SIZE),
				to_sfixed(-0.9846,1,L_SIZE),
				to_sfixed(-0.9846,1,L_SIZE),
				to_sfixed(-0.9846,1,L_SIZE),
				to_sfixed(-0.9846,1,L_SIZE),
				to_sfixed(-0.9846,1,L_SIZE),
				to_sfixed(-0.9845,1,L_SIZE),
				to_sfixed(-0.9845,1,L_SIZE),
				to_sfixed(-0.9845,1,L_SIZE),
				to_sfixed(-0.9845,1,L_SIZE),
				to_sfixed(-0.9845,1,L_SIZE),
				to_sfixed(-0.9845,1,L_SIZE),
				to_sfixed(-0.9845,1,L_SIZE),
				to_sfixed(-0.9845,1,L_SIZE),
				to_sfixed(-0.9845,1,L_SIZE),
				to_sfixed(-0.9844,1,L_SIZE),
				to_sfixed(-0.9844,1,L_SIZE),
				to_sfixed(-0.9844,1,L_SIZE),
				to_sfixed(-0.9844,1,L_SIZE),
				to_sfixed(-0.9844,1,L_SIZE),
				to_sfixed(-0.9844,1,L_SIZE),
				to_sfixed(-0.9844,1,L_SIZE),
				to_sfixed(-0.9844,1,L_SIZE),
				to_sfixed(-0.9844,1,L_SIZE),
				to_sfixed(-0.9843,1,L_SIZE),
				to_sfixed(-0.9843,1,L_SIZE),
				to_sfixed(-0.9843,1,L_SIZE),
				to_sfixed(-0.9843,1,L_SIZE),
				to_sfixed(-0.9843,1,L_SIZE),
				to_sfixed(-0.9843,1,L_SIZE),
				to_sfixed(-0.9843,1,L_SIZE),
				to_sfixed(-0.9843,1,L_SIZE),
				to_sfixed(-0.9843,1,L_SIZE),
				to_sfixed(-0.9842,1,L_SIZE),
				to_sfixed(-0.9842,1,L_SIZE),
				to_sfixed(-0.9842,1,L_SIZE),
				to_sfixed(-0.9842,1,L_SIZE),
				to_sfixed(-0.9842,1,L_SIZE),
				to_sfixed(-0.9842,1,L_SIZE),
				to_sfixed(-0.9842,1,L_SIZE),
				to_sfixed(-0.9842,1,L_SIZE),
				to_sfixed(-0.9841,1,L_SIZE),
				to_sfixed(-0.9841,1,L_SIZE),
				to_sfixed(-0.9841,1,L_SIZE),
				to_sfixed(-0.9841,1,L_SIZE),
				to_sfixed(-0.9841,1,L_SIZE),
				to_sfixed(-0.9841,1,L_SIZE),
				to_sfixed(-0.9841,1,L_SIZE),
				to_sfixed(-0.9841,1,L_SIZE),
				to_sfixed(-0.9841,1,L_SIZE),
				to_sfixed(-0.9840,1,L_SIZE),
				to_sfixed(-0.9840,1,L_SIZE),
				to_sfixed(-0.9840,1,L_SIZE),
				to_sfixed(-0.9840,1,L_SIZE),
				to_sfixed(-0.9840,1,L_SIZE),
				to_sfixed(-0.9840,1,L_SIZE),
				to_sfixed(-0.9840,1,L_SIZE),
				to_sfixed(-0.9840,1,L_SIZE),
				to_sfixed(-0.9840,1,L_SIZE),
				to_sfixed(-0.9839,1,L_SIZE),
				to_sfixed(-0.9839,1,L_SIZE),
				to_sfixed(-0.9839,1,L_SIZE),
				to_sfixed(-0.9839,1,L_SIZE),
				to_sfixed(-0.9839,1,L_SIZE),
				to_sfixed(-0.9839,1,L_SIZE),
				to_sfixed(-0.9839,1,L_SIZE),
				to_sfixed(-0.9839,1,L_SIZE),
				to_sfixed(-0.9838,1,L_SIZE),
				to_sfixed(-0.9838,1,L_SIZE),
				to_sfixed(-0.9838,1,L_SIZE),
				to_sfixed(-0.9838,1,L_SIZE),
				to_sfixed(-0.9838,1,L_SIZE),
				to_sfixed(-0.9838,1,L_SIZE),
				to_sfixed(-0.9838,1,L_SIZE),
				to_sfixed(-0.9838,1,L_SIZE),
				to_sfixed(-0.9838,1,L_SIZE),
				to_sfixed(-0.9837,1,L_SIZE),
				to_sfixed(-0.9837,1,L_SIZE),
				to_sfixed(-0.9837,1,L_SIZE),
				to_sfixed(-0.9837,1,L_SIZE),
				to_sfixed(-0.9837,1,L_SIZE),
				to_sfixed(-0.9837,1,L_SIZE),
				to_sfixed(-0.9837,1,L_SIZE),
				to_sfixed(-0.9837,1,L_SIZE),
				to_sfixed(-0.9836,1,L_SIZE),
				to_sfixed(-0.9836,1,L_SIZE),
				to_sfixed(-0.9836,1,L_SIZE),
				to_sfixed(-0.9836,1,L_SIZE),
				to_sfixed(-0.9836,1,L_SIZE),
				to_sfixed(-0.9836,1,L_SIZE),
				to_sfixed(-0.9836,1,L_SIZE),
				to_sfixed(-0.9836,1,L_SIZE),
				to_sfixed(-0.9835,1,L_SIZE),
				to_sfixed(-0.9835,1,L_SIZE),
				to_sfixed(-0.9835,1,L_SIZE),
				to_sfixed(-0.9835,1,L_SIZE),
				to_sfixed(-0.9835,1,L_SIZE),
				to_sfixed(-0.9835,1,L_SIZE),
				to_sfixed(-0.9835,1,L_SIZE),
				to_sfixed(-0.9835,1,L_SIZE),
				to_sfixed(-0.9835,1,L_SIZE),
				to_sfixed(-0.9834,1,L_SIZE),
				to_sfixed(-0.9834,1,L_SIZE),
				to_sfixed(-0.9834,1,L_SIZE),
				to_sfixed(-0.9834,1,L_SIZE),
				to_sfixed(-0.9834,1,L_SIZE),
				to_sfixed(-0.9834,1,L_SIZE),
				to_sfixed(-0.9834,1,L_SIZE),
				to_sfixed(-0.9834,1,L_SIZE),
				to_sfixed(-0.9833,1,L_SIZE),
				to_sfixed(-0.9833,1,L_SIZE),
				to_sfixed(-0.9833,1,L_SIZE),
				to_sfixed(-0.9833,1,L_SIZE),
				to_sfixed(-0.9833,1,L_SIZE),
				to_sfixed(-0.9833,1,L_SIZE),
				to_sfixed(-0.9833,1,L_SIZE),
				to_sfixed(-0.9833,1,L_SIZE),
				to_sfixed(-0.9832,1,L_SIZE),
				to_sfixed(-0.9832,1,L_SIZE),
				to_sfixed(-0.9832,1,L_SIZE),
				to_sfixed(-0.9832,1,L_SIZE),
				to_sfixed(-0.9832,1,L_SIZE),
				to_sfixed(-0.9832,1,L_SIZE),
				to_sfixed(-0.9832,1,L_SIZE),
				to_sfixed(-0.9832,1,L_SIZE),
				to_sfixed(-0.9831,1,L_SIZE),
				to_sfixed(-0.9831,1,L_SIZE),
				to_sfixed(-0.9831,1,L_SIZE),
				to_sfixed(-0.9831,1,L_SIZE),
				to_sfixed(-0.9831,1,L_SIZE),
				to_sfixed(-0.9831,1,L_SIZE),
				to_sfixed(-0.9831,1,L_SIZE),
				to_sfixed(-0.9831,1,L_SIZE),
				to_sfixed(-0.9831,1,L_SIZE),
				to_sfixed(-0.9830,1,L_SIZE),
				to_sfixed(-0.9830,1,L_SIZE),
				to_sfixed(-0.9830,1,L_SIZE),
				to_sfixed(-0.9830,1,L_SIZE),
				to_sfixed(-0.9830,1,L_SIZE),
				to_sfixed(-0.9830,1,L_SIZE),
				to_sfixed(-0.9830,1,L_SIZE),
				to_sfixed(-0.9830,1,L_SIZE),
				to_sfixed(-0.9829,1,L_SIZE),
				to_sfixed(-0.9829,1,L_SIZE),
				to_sfixed(-0.9829,1,L_SIZE),
				to_sfixed(-0.9829,1,L_SIZE),
				to_sfixed(-0.9829,1,L_SIZE),
				to_sfixed(-0.9829,1,L_SIZE),
				to_sfixed(-0.9829,1,L_SIZE),
				to_sfixed(-0.9829,1,L_SIZE),
				to_sfixed(-0.9828,1,L_SIZE),
				to_sfixed(-0.9828,1,L_SIZE),
				to_sfixed(-0.9828,1,L_SIZE),
				to_sfixed(-0.9828,1,L_SIZE),
				to_sfixed(-0.9828,1,L_SIZE),
				to_sfixed(-0.9828,1,L_SIZE),
				to_sfixed(-0.9828,1,L_SIZE),
				to_sfixed(-0.9828,1,L_SIZE),
				to_sfixed(-0.9827,1,L_SIZE),
				to_sfixed(-0.9827,1,L_SIZE),
				to_sfixed(-0.9827,1,L_SIZE),
				to_sfixed(-0.9827,1,L_SIZE),
				to_sfixed(-0.9827,1,L_SIZE),
				to_sfixed(-0.9827,1,L_SIZE),
				to_sfixed(-0.9827,1,L_SIZE),
				to_sfixed(-0.9827,1,L_SIZE),
				to_sfixed(-0.9826,1,L_SIZE),
				to_sfixed(-0.9826,1,L_SIZE),
				to_sfixed(-0.9826,1,L_SIZE),
				to_sfixed(-0.9826,1,L_SIZE),
				to_sfixed(-0.9826,1,L_SIZE),
				to_sfixed(-0.9826,1,L_SIZE),
				to_sfixed(-0.9826,1,L_SIZE),
				to_sfixed(-0.9826,1,L_SIZE),
				to_sfixed(-0.9825,1,L_SIZE),
				to_sfixed(-0.9825,1,L_SIZE),
				to_sfixed(-0.9825,1,L_SIZE),
				to_sfixed(-0.9825,1,L_SIZE),
				to_sfixed(-0.9825,1,L_SIZE),
				to_sfixed(-0.9825,1,L_SIZE),
				to_sfixed(-0.9825,1,L_SIZE),
				to_sfixed(-0.9825,1,L_SIZE),
				to_sfixed(-0.9824,1,L_SIZE),
				to_sfixed(-0.9824,1,L_SIZE),
				to_sfixed(-0.9824,1,L_SIZE),
				to_sfixed(-0.9824,1,L_SIZE),
				to_sfixed(-0.9824,1,L_SIZE),
				to_sfixed(-0.9824,1,L_SIZE),
				to_sfixed(-0.9824,1,L_SIZE),
				to_sfixed(-0.9823,1,L_SIZE),
				to_sfixed(-0.9823,1,L_SIZE),
				to_sfixed(-0.9823,1,L_SIZE),
				to_sfixed(-0.9823,1,L_SIZE),
				to_sfixed(-0.9823,1,L_SIZE),
				to_sfixed(-0.9823,1,L_SIZE),
				to_sfixed(-0.9823,1,L_SIZE),
				to_sfixed(-0.9823,1,L_SIZE),
				to_sfixed(-0.9822,1,L_SIZE),
				to_sfixed(-0.9822,1,L_SIZE),
				to_sfixed(-0.9822,1,L_SIZE),
				to_sfixed(-0.9822,1,L_SIZE),
				to_sfixed(-0.9822,1,L_SIZE),
				to_sfixed(-0.9822,1,L_SIZE),
				to_sfixed(-0.9822,1,L_SIZE),
				to_sfixed(-0.9822,1,L_SIZE),
				to_sfixed(-0.9821,1,L_SIZE),
				to_sfixed(-0.9821,1,L_SIZE),
				to_sfixed(-0.9821,1,L_SIZE),
				to_sfixed(-0.9821,1,L_SIZE),
				to_sfixed(-0.9821,1,L_SIZE),
				to_sfixed(-0.9821,1,L_SIZE),
				to_sfixed(-0.9821,1,L_SIZE),
				to_sfixed(-0.9821,1,L_SIZE),
				to_sfixed(-0.9820,1,L_SIZE),
				to_sfixed(-0.9820,1,L_SIZE),
				to_sfixed(-0.9820,1,L_SIZE),
				to_sfixed(-0.9820,1,L_SIZE),
				to_sfixed(-0.9820,1,L_SIZE),
				to_sfixed(-0.9820,1,L_SIZE),
				to_sfixed(-0.9820,1,L_SIZE),
				to_sfixed(-0.9819,1,L_SIZE),
				to_sfixed(-0.9819,1,L_SIZE),
				to_sfixed(-0.9819,1,L_SIZE),
				to_sfixed(-0.9819,1,L_SIZE),
				to_sfixed(-0.9819,1,L_SIZE),
				to_sfixed(-0.9819,1,L_SIZE),
				to_sfixed(-0.9819,1,L_SIZE),
				to_sfixed(-0.9819,1,L_SIZE),
				to_sfixed(-0.9818,1,L_SIZE),
				to_sfixed(-0.9818,1,L_SIZE),
				to_sfixed(-0.9818,1,L_SIZE),
				to_sfixed(-0.9818,1,L_SIZE),
				to_sfixed(-0.9818,1,L_SIZE),
				to_sfixed(-0.9818,1,L_SIZE),
				to_sfixed(-0.9818,1,L_SIZE),
				to_sfixed(-0.9817,1,L_SIZE),
				to_sfixed(-0.9817,1,L_SIZE),
				to_sfixed(-0.9817,1,L_SIZE),
				to_sfixed(-0.9817,1,L_SIZE),
				to_sfixed(-0.9817,1,L_SIZE),
				to_sfixed(-0.9817,1,L_SIZE),
				to_sfixed(-0.9817,1,L_SIZE),
				to_sfixed(-0.9817,1,L_SIZE),
				to_sfixed(-0.9816,1,L_SIZE),
				to_sfixed(-0.9816,1,L_SIZE),
				to_sfixed(-0.9816,1,L_SIZE),
				to_sfixed(-0.9816,1,L_SIZE),
				to_sfixed(-0.9816,1,L_SIZE),
				to_sfixed(-0.9816,1,L_SIZE),
				to_sfixed(-0.9816,1,L_SIZE),
				to_sfixed(-0.9815,1,L_SIZE),
				to_sfixed(-0.9815,1,L_SIZE),
				to_sfixed(-0.9815,1,L_SIZE),
				to_sfixed(-0.9815,1,L_SIZE),
				to_sfixed(-0.9815,1,L_SIZE),
				to_sfixed(-0.9815,1,L_SIZE),
				to_sfixed(-0.9815,1,L_SIZE),
				to_sfixed(-0.9815,1,L_SIZE),
				to_sfixed(-0.9814,1,L_SIZE),
				to_sfixed(-0.9814,1,L_SIZE),
				to_sfixed(-0.9814,1,L_SIZE),
				to_sfixed(-0.9814,1,L_SIZE),
				to_sfixed(-0.9814,1,L_SIZE),
				to_sfixed(-0.9814,1,L_SIZE),
				to_sfixed(-0.9814,1,L_SIZE),
				to_sfixed(-0.9813,1,L_SIZE),
				to_sfixed(-0.9813,1,L_SIZE),
				to_sfixed(-0.9813,1,L_SIZE),
				to_sfixed(-0.9813,1,L_SIZE),
				to_sfixed(-0.9813,1,L_SIZE),
				to_sfixed(-0.9813,1,L_SIZE),
				to_sfixed(-0.9813,1,L_SIZE),
				to_sfixed(-0.9813,1,L_SIZE),
				to_sfixed(-0.9812,1,L_SIZE),
				to_sfixed(-0.9812,1,L_SIZE),
				to_sfixed(-0.9812,1,L_SIZE),
				to_sfixed(-0.9812,1,L_SIZE),
				to_sfixed(-0.9812,1,L_SIZE),
				to_sfixed(-0.9812,1,L_SIZE),
				to_sfixed(-0.9812,1,L_SIZE),
				to_sfixed(-0.9811,1,L_SIZE),
				to_sfixed(-0.9811,1,L_SIZE),
				to_sfixed(-0.9811,1,L_SIZE),
				to_sfixed(-0.9811,1,L_SIZE),
				to_sfixed(-0.9811,1,L_SIZE),
				to_sfixed(-0.9811,1,L_SIZE),
				to_sfixed(-0.9811,1,L_SIZE),
				to_sfixed(-0.9810,1,L_SIZE),
				to_sfixed(-0.9810,1,L_SIZE),
				to_sfixed(-0.9810,1,L_SIZE),
				to_sfixed(-0.9810,1,L_SIZE),
				to_sfixed(-0.9810,1,L_SIZE),
				to_sfixed(-0.9810,1,L_SIZE),
				to_sfixed(-0.9810,1,L_SIZE),
				to_sfixed(-0.9810,1,L_SIZE),
				to_sfixed(-0.9809,1,L_SIZE),
				to_sfixed(-0.9809,1,L_SIZE),
				to_sfixed(-0.9809,1,L_SIZE),
				to_sfixed(-0.9809,1,L_SIZE),
				to_sfixed(-0.9809,1,L_SIZE),
				to_sfixed(-0.9809,1,L_SIZE),
				to_sfixed(-0.9809,1,L_SIZE),
				to_sfixed(-0.9808,1,L_SIZE),
				to_sfixed(-0.9808,1,L_SIZE),
				to_sfixed(-0.9808,1,L_SIZE),
				to_sfixed(-0.9808,1,L_SIZE),
				to_sfixed(-0.9808,1,L_SIZE),
				to_sfixed(-0.9808,1,L_SIZE),
				to_sfixed(-0.9808,1,L_SIZE),
				to_sfixed(-0.9807,1,L_SIZE),
				to_sfixed(-0.9807,1,L_SIZE),
				to_sfixed(-0.9807,1,L_SIZE),
				to_sfixed(-0.9807,1,L_SIZE),
				to_sfixed(-0.9807,1,L_SIZE),
				to_sfixed(-0.9807,1,L_SIZE),
				to_sfixed(-0.9807,1,L_SIZE),
				to_sfixed(-0.9806,1,L_SIZE),
				to_sfixed(-0.9806,1,L_SIZE),
				to_sfixed(-0.9806,1,L_SIZE),
				to_sfixed(-0.9806,1,L_SIZE),
				to_sfixed(-0.9806,1,L_SIZE),
				to_sfixed(-0.9806,1,L_SIZE),
				to_sfixed(-0.9806,1,L_SIZE),
				to_sfixed(-0.9805,1,L_SIZE),
				to_sfixed(-0.9805,1,L_SIZE),
				to_sfixed(-0.9805,1,L_SIZE),
				to_sfixed(-0.9805,1,L_SIZE),
				to_sfixed(-0.9805,1,L_SIZE),
				to_sfixed(-0.9805,1,L_SIZE),
				to_sfixed(-0.9805,1,L_SIZE),
				to_sfixed(-0.9804,1,L_SIZE),
				to_sfixed(-0.9804,1,L_SIZE),
				to_sfixed(-0.9804,1,L_SIZE),
				to_sfixed(-0.9804,1,L_SIZE),
				to_sfixed(-0.9804,1,L_SIZE),
				to_sfixed(-0.9804,1,L_SIZE),
				to_sfixed(-0.9804,1,L_SIZE),
				to_sfixed(-0.9803,1,L_SIZE),
				to_sfixed(-0.9803,1,L_SIZE),
				to_sfixed(-0.9803,1,L_SIZE),
				to_sfixed(-0.9803,1,L_SIZE),
				to_sfixed(-0.9803,1,L_SIZE),
				to_sfixed(-0.9803,1,L_SIZE),
				to_sfixed(-0.9803,1,L_SIZE),
				to_sfixed(-0.9802,1,L_SIZE),
				to_sfixed(-0.9802,1,L_SIZE),
				to_sfixed(-0.9802,1,L_SIZE),
				to_sfixed(-0.9802,1,L_SIZE),
				to_sfixed(-0.9802,1,L_SIZE),
				to_sfixed(-0.9802,1,L_SIZE),
				to_sfixed(-0.9802,1,L_SIZE),
				to_sfixed(-0.9801,1,L_SIZE),
				to_sfixed(-0.9801,1,L_SIZE),
				to_sfixed(-0.9801,1,L_SIZE),
				to_sfixed(-0.9801,1,L_SIZE),
				to_sfixed(-0.9801,1,L_SIZE),
				to_sfixed(-0.9801,1,L_SIZE),
				to_sfixed(-0.9801,1,L_SIZE),
				to_sfixed(-0.9800,1,L_SIZE),
				to_sfixed(-0.9800,1,L_SIZE),
				to_sfixed(-0.9800,1,L_SIZE),
				to_sfixed(-0.9800,1,L_SIZE),
				to_sfixed(-0.9800,1,L_SIZE),
				to_sfixed(-0.9800,1,L_SIZE),
				to_sfixed(-0.9800,1,L_SIZE),
				to_sfixed(-0.9799,1,L_SIZE),
				to_sfixed(-0.9799,1,L_SIZE),
				to_sfixed(-0.9799,1,L_SIZE),
				to_sfixed(-0.9799,1,L_SIZE),
				to_sfixed(-0.9799,1,L_SIZE),
				to_sfixed(-0.9799,1,L_SIZE),
				to_sfixed(-0.9799,1,L_SIZE),
				to_sfixed(-0.9798,1,L_SIZE),
				to_sfixed(-0.9798,1,L_SIZE),
				to_sfixed(-0.9798,1,L_SIZE),
				to_sfixed(-0.9798,1,L_SIZE),
				to_sfixed(-0.9798,1,L_SIZE),
				to_sfixed(-0.9798,1,L_SIZE),
				to_sfixed(-0.9798,1,L_SIZE),
				to_sfixed(-0.9797,1,L_SIZE),
				to_sfixed(-0.9797,1,L_SIZE),
				to_sfixed(-0.9797,1,L_SIZE),
				to_sfixed(-0.9797,1,L_SIZE),
				to_sfixed(-0.9797,1,L_SIZE),
				to_sfixed(-0.9797,1,L_SIZE),
				to_sfixed(-0.9797,1,L_SIZE),
				to_sfixed(-0.9796,1,L_SIZE),
				to_sfixed(-0.9796,1,L_SIZE),
				to_sfixed(-0.9796,1,L_SIZE),
				to_sfixed(-0.9796,1,L_SIZE),
				to_sfixed(-0.9796,1,L_SIZE),
				to_sfixed(-0.9796,1,L_SIZE),
				to_sfixed(-0.9795,1,L_SIZE),
				to_sfixed(-0.9795,1,L_SIZE),
				to_sfixed(-0.9795,1,L_SIZE),
				to_sfixed(-0.9795,1,L_SIZE),
				to_sfixed(-0.9795,1,L_SIZE),
				to_sfixed(-0.9795,1,L_SIZE),
				to_sfixed(-0.9795,1,L_SIZE),
				to_sfixed(-0.9794,1,L_SIZE),
				to_sfixed(-0.9794,1,L_SIZE),
				to_sfixed(-0.9794,1,L_SIZE),
				to_sfixed(-0.9794,1,L_SIZE),
				to_sfixed(-0.9794,1,L_SIZE),
				to_sfixed(-0.9794,1,L_SIZE),
				to_sfixed(-0.9794,1,L_SIZE),
				to_sfixed(-0.9793,1,L_SIZE),
				to_sfixed(-0.9793,1,L_SIZE),
				to_sfixed(-0.9793,1,L_SIZE),
				to_sfixed(-0.9793,1,L_SIZE),
				to_sfixed(-0.9793,1,L_SIZE),
				to_sfixed(-0.9793,1,L_SIZE),
				to_sfixed(-0.9792,1,L_SIZE),
				to_sfixed(-0.9792,1,L_SIZE),
				to_sfixed(-0.9792,1,L_SIZE),
				to_sfixed(-0.9792,1,L_SIZE),
				to_sfixed(-0.9792,1,L_SIZE),
				to_sfixed(-0.9792,1,L_SIZE),
				to_sfixed(-0.9792,1,L_SIZE),
				to_sfixed(-0.9791,1,L_SIZE),
				to_sfixed(-0.9791,1,L_SIZE),
				to_sfixed(-0.9791,1,L_SIZE),
				to_sfixed(-0.9791,1,L_SIZE),
				to_sfixed(-0.9791,1,L_SIZE),
				to_sfixed(-0.9791,1,L_SIZE),
				to_sfixed(-0.9791,1,L_SIZE),
				to_sfixed(-0.9790,1,L_SIZE),
				to_sfixed(-0.9790,1,L_SIZE),
				to_sfixed(-0.9790,1,L_SIZE),
				to_sfixed(-0.9790,1,L_SIZE),
				to_sfixed(-0.9790,1,L_SIZE),
				to_sfixed(-0.9790,1,L_SIZE),
				to_sfixed(-0.9789,1,L_SIZE),
				to_sfixed(-0.9789,1,L_SIZE),
				to_sfixed(-0.9789,1,L_SIZE),
				to_sfixed(-0.9789,1,L_SIZE),
				to_sfixed(-0.9789,1,L_SIZE),
				to_sfixed(-0.9789,1,L_SIZE),
				to_sfixed(-0.9789,1,L_SIZE),
				to_sfixed(-0.9788,1,L_SIZE),
				to_sfixed(-0.9788,1,L_SIZE),
				to_sfixed(-0.9788,1,L_SIZE),
				to_sfixed(-0.9788,1,L_SIZE),
				to_sfixed(-0.9788,1,L_SIZE),
				to_sfixed(-0.9788,1,L_SIZE),
				to_sfixed(-0.9787,1,L_SIZE),
				to_sfixed(-0.9787,1,L_SIZE),
				to_sfixed(-0.9787,1,L_SIZE),
				to_sfixed(-0.9787,1,L_SIZE),
				to_sfixed(-0.9787,1,L_SIZE),
				to_sfixed(-0.9787,1,L_SIZE),
				to_sfixed(-0.9787,1,L_SIZE),
				to_sfixed(-0.9786,1,L_SIZE),
				to_sfixed(-0.9786,1,L_SIZE),
				to_sfixed(-0.9786,1,L_SIZE),
				to_sfixed(-0.9786,1,L_SIZE),
				to_sfixed(-0.9786,1,L_SIZE),
				to_sfixed(-0.9786,1,L_SIZE),
				to_sfixed(-0.9785,1,L_SIZE),
				to_sfixed(-0.9785,1,L_SIZE),
				to_sfixed(-0.9785,1,L_SIZE),
				to_sfixed(-0.9785,1,L_SIZE),
				to_sfixed(-0.9785,1,L_SIZE),
				to_sfixed(-0.9785,1,L_SIZE),
				to_sfixed(-0.9785,1,L_SIZE),
				to_sfixed(-0.9784,1,L_SIZE),
				to_sfixed(-0.9784,1,L_SIZE),
				to_sfixed(-0.9784,1,L_SIZE),
				to_sfixed(-0.9784,1,L_SIZE),
				to_sfixed(-0.9784,1,L_SIZE),
				to_sfixed(-0.9784,1,L_SIZE),
				to_sfixed(-0.9783,1,L_SIZE),
				to_sfixed(-0.9783,1,L_SIZE),
				to_sfixed(-0.9783,1,L_SIZE),
				to_sfixed(-0.9783,1,L_SIZE),
				to_sfixed(-0.9783,1,L_SIZE),
				to_sfixed(-0.9783,1,L_SIZE),
				to_sfixed(-0.9782,1,L_SIZE),
				to_sfixed(-0.9782,1,L_SIZE),
				to_sfixed(-0.9782,1,L_SIZE),
				to_sfixed(-0.9782,1,L_SIZE),
				to_sfixed(-0.9782,1,L_SIZE),
				to_sfixed(-0.9782,1,L_SIZE),
				to_sfixed(-0.9782,1,L_SIZE),
				to_sfixed(-0.9781,1,L_SIZE),
				to_sfixed(-0.9781,1,L_SIZE),
				to_sfixed(-0.9781,1,L_SIZE),
				to_sfixed(-0.9781,1,L_SIZE),
				to_sfixed(-0.9781,1,L_SIZE),
				to_sfixed(-0.9781,1,L_SIZE),
				to_sfixed(-0.9780,1,L_SIZE),
				to_sfixed(-0.9780,1,L_SIZE),
				to_sfixed(-0.9780,1,L_SIZE),
				to_sfixed(-0.9780,1,L_SIZE),
				to_sfixed(-0.9780,1,L_SIZE),
				to_sfixed(-0.9780,1,L_SIZE),
				to_sfixed(-0.9779,1,L_SIZE),
				to_sfixed(-0.9779,1,L_SIZE),
				to_sfixed(-0.9779,1,L_SIZE),
				to_sfixed(-0.9779,1,L_SIZE),
				to_sfixed(-0.9779,1,L_SIZE),
				to_sfixed(-0.9779,1,L_SIZE),
				to_sfixed(-0.9779,1,L_SIZE),
				to_sfixed(-0.9778,1,L_SIZE),
				to_sfixed(-0.9778,1,L_SIZE),
				to_sfixed(-0.9778,1,L_SIZE),
				to_sfixed(-0.9778,1,L_SIZE),
				to_sfixed(-0.9778,1,L_SIZE),
				to_sfixed(-0.9778,1,L_SIZE),
				to_sfixed(-0.9777,1,L_SIZE),
				to_sfixed(-0.9777,1,L_SIZE),
				to_sfixed(-0.9777,1,L_SIZE),
				to_sfixed(-0.9777,1,L_SIZE),
				to_sfixed(-0.9777,1,L_SIZE),
				to_sfixed(-0.9777,1,L_SIZE),
				to_sfixed(-0.9776,1,L_SIZE),
				to_sfixed(-0.9776,1,L_SIZE),
				to_sfixed(-0.9776,1,L_SIZE),
				to_sfixed(-0.9776,1,L_SIZE),
				to_sfixed(-0.9776,1,L_SIZE),
				to_sfixed(-0.9776,1,L_SIZE),
				to_sfixed(-0.9775,1,L_SIZE),
				to_sfixed(-0.9775,1,L_SIZE),
				to_sfixed(-0.9775,1,L_SIZE),
				to_sfixed(-0.9775,1,L_SIZE),
				to_sfixed(-0.9775,1,L_SIZE),
				to_sfixed(-0.9775,1,L_SIZE),
				to_sfixed(-0.9774,1,L_SIZE),
				to_sfixed(-0.9774,1,L_SIZE),
				to_sfixed(-0.9774,1,L_SIZE),
				to_sfixed(-0.9774,1,L_SIZE),
				to_sfixed(-0.9774,1,L_SIZE),
				to_sfixed(-0.9774,1,L_SIZE),
				to_sfixed(-0.9773,1,L_SIZE),
				to_sfixed(-0.9773,1,L_SIZE),
				to_sfixed(-0.9773,1,L_SIZE),
				to_sfixed(-0.9773,1,L_SIZE),
				to_sfixed(-0.9773,1,L_SIZE),
				to_sfixed(-0.9773,1,L_SIZE),
				to_sfixed(-0.9772,1,L_SIZE),
				to_sfixed(-0.9772,1,L_SIZE),
				to_sfixed(-0.9772,1,L_SIZE),
				to_sfixed(-0.9772,1,L_SIZE),
				to_sfixed(-0.9772,1,L_SIZE),
				to_sfixed(-0.9772,1,L_SIZE),
				to_sfixed(-0.9771,1,L_SIZE),
				to_sfixed(-0.9771,1,L_SIZE),
				to_sfixed(-0.9771,1,L_SIZE),
				to_sfixed(-0.9771,1,L_SIZE),
				to_sfixed(-0.9771,1,L_SIZE),
				to_sfixed(-0.9771,1,L_SIZE),
				to_sfixed(-0.9771,1,L_SIZE),
				to_sfixed(-0.9770,1,L_SIZE),
				to_sfixed(-0.9770,1,L_SIZE),
				to_sfixed(-0.9770,1,L_SIZE),
				to_sfixed(-0.9770,1,L_SIZE),
				to_sfixed(-0.9770,1,L_SIZE),
				to_sfixed(-0.9770,1,L_SIZE),
				to_sfixed(-0.9769,1,L_SIZE),
				to_sfixed(-0.9769,1,L_SIZE),
				to_sfixed(-0.9769,1,L_SIZE),
				to_sfixed(-0.9769,1,L_SIZE),
				to_sfixed(-0.9769,1,L_SIZE),
				to_sfixed(-0.9769,1,L_SIZE),
				to_sfixed(-0.9768,1,L_SIZE),
				to_sfixed(-0.9768,1,L_SIZE),
				to_sfixed(-0.9768,1,L_SIZE),
				to_sfixed(-0.9768,1,L_SIZE),
				to_sfixed(-0.9768,1,L_SIZE),
				to_sfixed(-0.9767,1,L_SIZE),
				to_sfixed(-0.9767,1,L_SIZE),
				to_sfixed(-0.9767,1,L_SIZE),
				to_sfixed(-0.9767,1,L_SIZE),
				to_sfixed(-0.9767,1,L_SIZE),
				to_sfixed(-0.9767,1,L_SIZE),
				to_sfixed(-0.9766,1,L_SIZE),
				to_sfixed(-0.9766,1,L_SIZE),
				to_sfixed(-0.9766,1,L_SIZE),
				to_sfixed(-0.9766,1,L_SIZE),
				to_sfixed(-0.9766,1,L_SIZE),
				to_sfixed(-0.9766,1,L_SIZE),
				to_sfixed(-0.9765,1,L_SIZE),
				to_sfixed(-0.9765,1,L_SIZE),
				to_sfixed(-0.9765,1,L_SIZE),
				to_sfixed(-0.9765,1,L_SIZE),
				to_sfixed(-0.9765,1,L_SIZE),
				to_sfixed(-0.9765,1,L_SIZE),
				to_sfixed(-0.9764,1,L_SIZE),
				to_sfixed(-0.9764,1,L_SIZE),
				to_sfixed(-0.9764,1,L_SIZE),
				to_sfixed(-0.9764,1,L_SIZE),
				to_sfixed(-0.9764,1,L_SIZE),
				to_sfixed(-0.9764,1,L_SIZE),
				to_sfixed(-0.9763,1,L_SIZE),
				to_sfixed(-0.9763,1,L_SIZE),
				to_sfixed(-0.9763,1,L_SIZE),
				to_sfixed(-0.9763,1,L_SIZE),
				to_sfixed(-0.9763,1,L_SIZE),
				to_sfixed(-0.9763,1,L_SIZE),
				to_sfixed(-0.9762,1,L_SIZE),
				to_sfixed(-0.9762,1,L_SIZE),
				to_sfixed(-0.9762,1,L_SIZE),
				to_sfixed(-0.9762,1,L_SIZE),
				to_sfixed(-0.9762,1,L_SIZE),
				to_sfixed(-0.9762,1,L_SIZE),
				to_sfixed(-0.9761,1,L_SIZE),
				to_sfixed(-0.9761,1,L_SIZE),
				to_sfixed(-0.9761,1,L_SIZE),
				to_sfixed(-0.9761,1,L_SIZE),
				to_sfixed(-0.9761,1,L_SIZE),
				to_sfixed(-0.9760,1,L_SIZE),
				to_sfixed(-0.9760,1,L_SIZE),
				to_sfixed(-0.9760,1,L_SIZE),
				to_sfixed(-0.9760,1,L_SIZE),
				to_sfixed(-0.9760,1,L_SIZE),
				to_sfixed(-0.9760,1,L_SIZE),
				to_sfixed(-0.9759,1,L_SIZE),
				to_sfixed(-0.9759,1,L_SIZE),
				to_sfixed(-0.9759,1,L_SIZE),
				to_sfixed(-0.9759,1,L_SIZE),
				to_sfixed(-0.9759,1,L_SIZE),
				to_sfixed(-0.9759,1,L_SIZE),
				to_sfixed(-0.9758,1,L_SIZE),
				to_sfixed(-0.9758,1,L_SIZE),
				to_sfixed(-0.9758,1,L_SIZE),
				to_sfixed(-0.9758,1,L_SIZE),
				to_sfixed(-0.9758,1,L_SIZE),
				to_sfixed(-0.9758,1,L_SIZE),
				to_sfixed(-0.9757,1,L_SIZE),
				to_sfixed(-0.9757,1,L_SIZE),
				to_sfixed(-0.9757,1,L_SIZE),
				to_sfixed(-0.9757,1,L_SIZE),
				to_sfixed(-0.9757,1,L_SIZE),
				to_sfixed(-0.9756,1,L_SIZE),
				to_sfixed(-0.9756,1,L_SIZE),
				to_sfixed(-0.9756,1,L_SIZE),
				to_sfixed(-0.9756,1,L_SIZE),
				to_sfixed(-0.9756,1,L_SIZE),
				to_sfixed(-0.9756,1,L_SIZE),
				to_sfixed(-0.9755,1,L_SIZE),
				to_sfixed(-0.9755,1,L_SIZE),
				to_sfixed(-0.9755,1,L_SIZE),
				to_sfixed(-0.9755,1,L_SIZE),
				to_sfixed(-0.9755,1,L_SIZE),
				to_sfixed(-0.9755,1,L_SIZE),
				to_sfixed(-0.9754,1,L_SIZE),
				to_sfixed(-0.9754,1,L_SIZE),
				to_sfixed(-0.9754,1,L_SIZE),
				to_sfixed(-0.9754,1,L_SIZE),
				to_sfixed(-0.9754,1,L_SIZE),
				to_sfixed(-0.9753,1,L_SIZE),
				to_sfixed(-0.9753,1,L_SIZE),
				to_sfixed(-0.9753,1,L_SIZE),
				to_sfixed(-0.9753,1,L_SIZE),
				to_sfixed(-0.9753,1,L_SIZE),
				to_sfixed(-0.9753,1,L_SIZE),
				to_sfixed(-0.9752,1,L_SIZE),
				to_sfixed(-0.9752,1,L_SIZE),
				to_sfixed(-0.9752,1,L_SIZE),
				to_sfixed(-0.9752,1,L_SIZE),
				to_sfixed(-0.9752,1,L_SIZE),
				to_sfixed(-0.9751,1,L_SIZE),
				to_sfixed(-0.9751,1,L_SIZE),
				to_sfixed(-0.9751,1,L_SIZE),
				to_sfixed(-0.9751,1,L_SIZE),
				to_sfixed(-0.9751,1,L_SIZE),
				to_sfixed(-0.9751,1,L_SIZE),
				to_sfixed(-0.9750,1,L_SIZE),
				to_sfixed(-0.9750,1,L_SIZE),
				to_sfixed(-0.9750,1,L_SIZE),
				to_sfixed(-0.9750,1,L_SIZE),
				to_sfixed(-0.9750,1,L_SIZE),
				to_sfixed(-0.9750,1,L_SIZE),
				to_sfixed(-0.9749,1,L_SIZE),
				to_sfixed(-0.9749,1,L_SIZE),
				to_sfixed(-0.9749,1,L_SIZE),
				to_sfixed(-0.9749,1,L_SIZE),
				to_sfixed(-0.9749,1,L_SIZE),
				to_sfixed(-0.9748,1,L_SIZE),
				to_sfixed(-0.9748,1,L_SIZE),
				to_sfixed(-0.9748,1,L_SIZE),
				to_sfixed(-0.9748,1,L_SIZE),
				to_sfixed(-0.9748,1,L_SIZE),
				to_sfixed(-0.9748,1,L_SIZE),
				to_sfixed(-0.9747,1,L_SIZE),
				to_sfixed(-0.9747,1,L_SIZE),
				to_sfixed(-0.9747,1,L_SIZE),
				to_sfixed(-0.9747,1,L_SIZE),
				to_sfixed(-0.9747,1,L_SIZE),
				to_sfixed(-0.9746,1,L_SIZE),
				to_sfixed(-0.9746,1,L_SIZE),
				to_sfixed(-0.9746,1,L_SIZE),
				to_sfixed(-0.9746,1,L_SIZE),
				to_sfixed(-0.9746,1,L_SIZE),
				to_sfixed(-0.9745,1,L_SIZE),
				to_sfixed(-0.9745,1,L_SIZE),
				to_sfixed(-0.9745,1,L_SIZE),
				to_sfixed(-0.9745,1,L_SIZE),
				to_sfixed(-0.9745,1,L_SIZE),
				to_sfixed(-0.9745,1,L_SIZE),
				to_sfixed(-0.9744,1,L_SIZE),
				to_sfixed(-0.9744,1,L_SIZE),
				to_sfixed(-0.9744,1,L_SIZE),
				to_sfixed(-0.9744,1,L_SIZE),
				to_sfixed(-0.9744,1,L_SIZE),
				to_sfixed(-0.9743,1,L_SIZE),
				to_sfixed(-0.9743,1,L_SIZE),
				to_sfixed(-0.9743,1,L_SIZE),
				to_sfixed(-0.9743,1,L_SIZE),
				to_sfixed(-0.9743,1,L_SIZE),
				to_sfixed(-0.9743,1,L_SIZE),
				to_sfixed(-0.9742,1,L_SIZE),
				to_sfixed(-0.9742,1,L_SIZE),
				to_sfixed(-0.9742,1,L_SIZE),
				to_sfixed(-0.9742,1,L_SIZE),
				to_sfixed(-0.9742,1,L_SIZE),
				to_sfixed(-0.9741,1,L_SIZE),
				to_sfixed(-0.9741,1,L_SIZE),
				to_sfixed(-0.9741,1,L_SIZE),
				to_sfixed(-0.9741,1,L_SIZE),
				to_sfixed(-0.9741,1,L_SIZE),
				to_sfixed(-0.9740,1,L_SIZE),
				to_sfixed(-0.9740,1,L_SIZE),
				to_sfixed(-0.9740,1,L_SIZE),
				to_sfixed(-0.9740,1,L_SIZE),
				to_sfixed(-0.9740,1,L_SIZE),
				to_sfixed(-0.9740,1,L_SIZE),
				to_sfixed(-0.9739,1,L_SIZE),
				to_sfixed(-0.9739,1,L_SIZE),
				to_sfixed(-0.9739,1,L_SIZE),
				to_sfixed(-0.9739,1,L_SIZE),
				to_sfixed(-0.9739,1,L_SIZE),
				to_sfixed(-0.9738,1,L_SIZE),
				to_sfixed(-0.9738,1,L_SIZE),
				to_sfixed(-0.9738,1,L_SIZE),
				to_sfixed(-0.9738,1,L_SIZE),
				to_sfixed(-0.9738,1,L_SIZE),
				to_sfixed(-0.9737,1,L_SIZE),
				to_sfixed(-0.9737,1,L_SIZE),
				to_sfixed(-0.9737,1,L_SIZE),
				to_sfixed(-0.9737,1,L_SIZE),
				to_sfixed(-0.9737,1,L_SIZE),
				to_sfixed(-0.9736,1,L_SIZE),
				to_sfixed(-0.9736,1,L_SIZE),
				to_sfixed(-0.9736,1,L_SIZE),
				to_sfixed(-0.9736,1,L_SIZE),
				to_sfixed(-0.9736,1,L_SIZE),
				to_sfixed(-0.9736,1,L_SIZE),
				to_sfixed(-0.9735,1,L_SIZE),
				to_sfixed(-0.9735,1,L_SIZE),
				to_sfixed(-0.9735,1,L_SIZE),
				to_sfixed(-0.9735,1,L_SIZE),
				to_sfixed(-0.9735,1,L_SIZE),
				to_sfixed(-0.9734,1,L_SIZE),
				to_sfixed(-0.9734,1,L_SIZE),
				to_sfixed(-0.9734,1,L_SIZE),
				to_sfixed(-0.9734,1,L_SIZE),
				to_sfixed(-0.9734,1,L_SIZE),
				to_sfixed(-0.9733,1,L_SIZE),
				to_sfixed(-0.9733,1,L_SIZE),
				to_sfixed(-0.9733,1,L_SIZE),
				to_sfixed(-0.9733,1,L_SIZE),
				to_sfixed(-0.9733,1,L_SIZE),
				to_sfixed(-0.9732,1,L_SIZE),
				to_sfixed(-0.9732,1,L_SIZE),
				to_sfixed(-0.9732,1,L_SIZE),
				to_sfixed(-0.9732,1,L_SIZE),
				to_sfixed(-0.9732,1,L_SIZE),
				to_sfixed(-0.9731,1,L_SIZE),
				to_sfixed(-0.9731,1,L_SIZE),
				to_sfixed(-0.9731,1,L_SIZE),
				to_sfixed(-0.9731,1,L_SIZE),
				to_sfixed(-0.9731,1,L_SIZE),
				to_sfixed(-0.9731,1,L_SIZE),
				to_sfixed(-0.9730,1,L_SIZE),
				to_sfixed(-0.9730,1,L_SIZE),
				to_sfixed(-0.9730,1,L_SIZE),
				to_sfixed(-0.9730,1,L_SIZE),
				to_sfixed(-0.9730,1,L_SIZE),
				to_sfixed(-0.9729,1,L_SIZE),
				to_sfixed(-0.9729,1,L_SIZE),
				to_sfixed(-0.9729,1,L_SIZE),
				to_sfixed(-0.9729,1,L_SIZE),
				to_sfixed(-0.9729,1,L_SIZE),
				to_sfixed(-0.9728,1,L_SIZE),
				to_sfixed(-0.9728,1,L_SIZE),
				to_sfixed(-0.9728,1,L_SIZE),
				to_sfixed(-0.9728,1,L_SIZE),
				to_sfixed(-0.9728,1,L_SIZE),
				to_sfixed(-0.9727,1,L_SIZE),
				to_sfixed(-0.9727,1,L_SIZE),
				to_sfixed(-0.9727,1,L_SIZE),
				to_sfixed(-0.9727,1,L_SIZE),
				to_sfixed(-0.9727,1,L_SIZE),
				to_sfixed(-0.9726,1,L_SIZE),
				to_sfixed(-0.9726,1,L_SIZE),
				to_sfixed(-0.9726,1,L_SIZE),
				to_sfixed(-0.9726,1,L_SIZE),
				to_sfixed(-0.9726,1,L_SIZE),
				to_sfixed(-0.9725,1,L_SIZE),
				to_sfixed(-0.9725,1,L_SIZE),
				to_sfixed(-0.9725,1,L_SIZE),
				to_sfixed(-0.9725,1,L_SIZE),
				to_sfixed(-0.9725,1,L_SIZE),
				to_sfixed(-0.9724,1,L_SIZE),
				to_sfixed(-0.9724,1,L_SIZE),
				to_sfixed(-0.9724,1,L_SIZE),
				to_sfixed(-0.9724,1,L_SIZE),
				to_sfixed(-0.9724,1,L_SIZE),
				to_sfixed(-0.9723,1,L_SIZE),
				to_sfixed(-0.9723,1,L_SIZE),
				to_sfixed(-0.9723,1,L_SIZE),
				to_sfixed(-0.9723,1,L_SIZE),
				to_sfixed(-0.9723,1,L_SIZE),
				to_sfixed(-0.9722,1,L_SIZE),
				to_sfixed(-0.9722,1,L_SIZE),
				to_sfixed(-0.9722,1,L_SIZE),
				to_sfixed(-0.9722,1,L_SIZE),
				to_sfixed(-0.9722,1,L_SIZE),
				to_sfixed(-0.9721,1,L_SIZE),
				to_sfixed(-0.9721,1,L_SIZE),
				to_sfixed(-0.9721,1,L_SIZE),
				to_sfixed(-0.9721,1,L_SIZE),
				to_sfixed(-0.9721,1,L_SIZE),
				to_sfixed(-0.9720,1,L_SIZE),
				to_sfixed(-0.9720,1,L_SIZE),
				to_sfixed(-0.9720,1,L_SIZE),
				to_sfixed(-0.9720,1,L_SIZE),
				to_sfixed(-0.9720,1,L_SIZE),
				to_sfixed(-0.9719,1,L_SIZE),
				to_sfixed(-0.9719,1,L_SIZE),
				to_sfixed(-0.9719,1,L_SIZE),
				to_sfixed(-0.9719,1,L_SIZE),
				to_sfixed(-0.9719,1,L_SIZE),
				to_sfixed(-0.9718,1,L_SIZE),
				to_sfixed(-0.9718,1,L_SIZE),
				to_sfixed(-0.9718,1,L_SIZE),
				to_sfixed(-0.9718,1,L_SIZE),
				to_sfixed(-0.9718,1,L_SIZE),
				to_sfixed(-0.9717,1,L_SIZE),
				to_sfixed(-0.9717,1,L_SIZE),
				to_sfixed(-0.9717,1,L_SIZE),
				to_sfixed(-0.9717,1,L_SIZE),
				to_sfixed(-0.9717,1,L_SIZE),
				to_sfixed(-0.9716,1,L_SIZE),
				to_sfixed(-0.9716,1,L_SIZE),
				to_sfixed(-0.9716,1,L_SIZE),
				to_sfixed(-0.9716,1,L_SIZE),
				to_sfixed(-0.9716,1,L_SIZE),
				to_sfixed(-0.9715,1,L_SIZE),
				to_sfixed(-0.9715,1,L_SIZE),
				to_sfixed(-0.9715,1,L_SIZE),
				to_sfixed(-0.9715,1,L_SIZE),
				to_sfixed(-0.9714,1,L_SIZE),
				to_sfixed(-0.9714,1,L_SIZE),
				to_sfixed(-0.9714,1,L_SIZE),
				to_sfixed(-0.9714,1,L_SIZE),
				to_sfixed(-0.9714,1,L_SIZE),
				to_sfixed(-0.9713,1,L_SIZE),
				to_sfixed(-0.9713,1,L_SIZE),
				to_sfixed(-0.9713,1,L_SIZE),
				to_sfixed(-0.9713,1,L_SIZE),
				to_sfixed(-0.9713,1,L_SIZE),
				to_sfixed(-0.9712,1,L_SIZE),
				to_sfixed(-0.9712,1,L_SIZE),
				to_sfixed(-0.9712,1,L_SIZE),
				to_sfixed(-0.9712,1,L_SIZE),
				to_sfixed(-0.9712,1,L_SIZE),
				to_sfixed(-0.9711,1,L_SIZE),
				to_sfixed(-0.9711,1,L_SIZE),
				to_sfixed(-0.9711,1,L_SIZE),
				to_sfixed(-0.9711,1,L_SIZE),
				to_sfixed(-0.9711,1,L_SIZE),
				to_sfixed(-0.9710,1,L_SIZE),
				to_sfixed(-0.9710,1,L_SIZE),
				to_sfixed(-0.9710,1,L_SIZE),
				to_sfixed(-0.9710,1,L_SIZE),
				to_sfixed(-0.9710,1,L_SIZE),
				to_sfixed(-0.9709,1,L_SIZE),
				to_sfixed(-0.9709,1,L_SIZE),
				to_sfixed(-0.9709,1,L_SIZE),
				to_sfixed(-0.9709,1,L_SIZE),
				to_sfixed(-0.9708,1,L_SIZE),
				to_sfixed(-0.9708,1,L_SIZE),
				to_sfixed(-0.9708,1,L_SIZE),
				to_sfixed(-0.9708,1,L_SIZE),
				to_sfixed(-0.9708,1,L_SIZE),
				to_sfixed(-0.9707,1,L_SIZE),
				to_sfixed(-0.9707,1,L_SIZE),
				to_sfixed(-0.9707,1,L_SIZE),
				to_sfixed(-0.9707,1,L_SIZE),
				to_sfixed(-0.9707,1,L_SIZE),
				to_sfixed(-0.9706,1,L_SIZE),
				to_sfixed(-0.9706,1,L_SIZE),
				to_sfixed(-0.9706,1,L_SIZE),
				to_sfixed(-0.9706,1,L_SIZE),
				to_sfixed(-0.9705,1,L_SIZE),
				to_sfixed(-0.9705,1,L_SIZE),
				to_sfixed(-0.9705,1,L_SIZE),
				to_sfixed(-0.9705,1,L_SIZE),
				to_sfixed(-0.9705,1,L_SIZE),
				to_sfixed(-0.9704,1,L_SIZE),
				to_sfixed(-0.9704,1,L_SIZE),
				to_sfixed(-0.9704,1,L_SIZE),
				to_sfixed(-0.9704,1,L_SIZE),
				to_sfixed(-0.9704,1,L_SIZE),
				to_sfixed(-0.9703,1,L_SIZE),
				to_sfixed(-0.9703,1,L_SIZE),
				to_sfixed(-0.9703,1,L_SIZE),
				to_sfixed(-0.9703,1,L_SIZE),
				to_sfixed(-0.9703,1,L_SIZE),
				to_sfixed(-0.9702,1,L_SIZE),
				to_sfixed(-0.9702,1,L_SIZE),
				to_sfixed(-0.9702,1,L_SIZE),
				to_sfixed(-0.9702,1,L_SIZE),
				to_sfixed(-0.9701,1,L_SIZE),
				to_sfixed(-0.9701,1,L_SIZE),
				to_sfixed(-0.9701,1,L_SIZE),
				to_sfixed(-0.9701,1,L_SIZE),
				to_sfixed(-0.9701,1,L_SIZE),
				to_sfixed(-0.9700,1,L_SIZE),
				to_sfixed(-0.9700,1,L_SIZE),
				to_sfixed(-0.9700,1,L_SIZE),
				to_sfixed(-0.9700,1,L_SIZE),
				to_sfixed(-0.9699,1,L_SIZE),
				to_sfixed(-0.9699,1,L_SIZE),
				to_sfixed(-0.9699,1,L_SIZE),
				to_sfixed(-0.9699,1,L_SIZE),
				to_sfixed(-0.9699,1,L_SIZE),
				to_sfixed(-0.9698,1,L_SIZE),
				to_sfixed(-0.9698,1,L_SIZE),
				to_sfixed(-0.9698,1,L_SIZE),
				to_sfixed(-0.9698,1,L_SIZE),
				to_sfixed(-0.9698,1,L_SIZE),
				to_sfixed(-0.9697,1,L_SIZE),
				to_sfixed(-0.9697,1,L_SIZE),
				to_sfixed(-0.9697,1,L_SIZE),
				to_sfixed(-0.9697,1,L_SIZE),
				to_sfixed(-0.9696,1,L_SIZE),
				to_sfixed(-0.9696,1,L_SIZE),
				to_sfixed(-0.9696,1,L_SIZE),
				to_sfixed(-0.9696,1,L_SIZE),
				to_sfixed(-0.9696,1,L_SIZE),
				to_sfixed(-0.9695,1,L_SIZE),
				to_sfixed(-0.9695,1,L_SIZE),
				to_sfixed(-0.9695,1,L_SIZE),
				to_sfixed(-0.9695,1,L_SIZE),
				to_sfixed(-0.9694,1,L_SIZE),
				to_sfixed(-0.9694,1,L_SIZE),
				to_sfixed(-0.9694,1,L_SIZE),
				to_sfixed(-0.9694,1,L_SIZE),
				to_sfixed(-0.9694,1,L_SIZE),
				to_sfixed(-0.9693,1,L_SIZE),
				to_sfixed(-0.9693,1,L_SIZE),
				to_sfixed(-0.9693,1,L_SIZE),
				to_sfixed(-0.9693,1,L_SIZE),
				to_sfixed(-0.9692,1,L_SIZE),
				to_sfixed(-0.9692,1,L_SIZE),
				to_sfixed(-0.9692,1,L_SIZE),
				to_sfixed(-0.9692,1,L_SIZE),
				to_sfixed(-0.9692,1,L_SIZE),
				to_sfixed(-0.9691,1,L_SIZE),
				to_sfixed(-0.9691,1,L_SIZE),
				to_sfixed(-0.9691,1,L_SIZE),
				to_sfixed(-0.9691,1,L_SIZE),
				to_sfixed(-0.9690,1,L_SIZE),
				to_sfixed(-0.9690,1,L_SIZE),
				to_sfixed(-0.9690,1,L_SIZE),
				to_sfixed(-0.9690,1,L_SIZE),
				to_sfixed(-0.9690,1,L_SIZE),
				to_sfixed(-0.9689,1,L_SIZE),
				to_sfixed(-0.9689,1,L_SIZE),
				to_sfixed(-0.9689,1,L_SIZE),
				to_sfixed(-0.9689,1,L_SIZE),
				to_sfixed(-0.9688,1,L_SIZE),
				to_sfixed(-0.9688,1,L_SIZE),
				to_sfixed(-0.9688,1,L_SIZE),
				to_sfixed(-0.9688,1,L_SIZE),
				to_sfixed(-0.9688,1,L_SIZE),
				to_sfixed(-0.9687,1,L_SIZE),
				to_sfixed(-0.9687,1,L_SIZE),
				to_sfixed(-0.9687,1,L_SIZE),
				to_sfixed(-0.9687,1,L_SIZE),
				to_sfixed(-0.9686,1,L_SIZE),
				to_sfixed(-0.9686,1,L_SIZE),
				to_sfixed(-0.9686,1,L_SIZE),
				to_sfixed(-0.9686,1,L_SIZE),
				to_sfixed(-0.9686,1,L_SIZE),
				to_sfixed(-0.9685,1,L_SIZE),
				to_sfixed(-0.9685,1,L_SIZE),
				to_sfixed(-0.9685,1,L_SIZE),
				to_sfixed(-0.9685,1,L_SIZE),
				to_sfixed(-0.9684,1,L_SIZE),
				to_sfixed(-0.9684,1,L_SIZE),
				to_sfixed(-0.9684,1,L_SIZE),
				to_sfixed(-0.9684,1,L_SIZE),
				to_sfixed(-0.9683,1,L_SIZE),
				to_sfixed(-0.9683,1,L_SIZE),
				to_sfixed(-0.9683,1,L_SIZE),
				to_sfixed(-0.9683,1,L_SIZE),
				to_sfixed(-0.9683,1,L_SIZE),
				to_sfixed(-0.9682,1,L_SIZE),
				to_sfixed(-0.9682,1,L_SIZE),
				to_sfixed(-0.9682,1,L_SIZE),
				to_sfixed(-0.9682,1,L_SIZE),
				to_sfixed(-0.9681,1,L_SIZE),
				to_sfixed(-0.9681,1,L_SIZE),
				to_sfixed(-0.9681,1,L_SIZE),
				to_sfixed(-0.9681,1,L_SIZE),
				to_sfixed(-0.9680,1,L_SIZE),
				to_sfixed(-0.9680,1,L_SIZE),
				to_sfixed(-0.9680,1,L_SIZE),
				to_sfixed(-0.9680,1,L_SIZE),
				to_sfixed(-0.9680,1,L_SIZE),
				to_sfixed(-0.9679,1,L_SIZE),
				to_sfixed(-0.9679,1,L_SIZE),
				to_sfixed(-0.9679,1,L_SIZE),
				to_sfixed(-0.9679,1,L_SIZE),
				to_sfixed(-0.9678,1,L_SIZE),
				to_sfixed(-0.9678,1,L_SIZE),
				to_sfixed(-0.9678,1,L_SIZE),
				to_sfixed(-0.9678,1,L_SIZE),
				to_sfixed(-0.9677,1,L_SIZE),
				to_sfixed(-0.9677,1,L_SIZE),
				to_sfixed(-0.9677,1,L_SIZE),
				to_sfixed(-0.9677,1,L_SIZE),
				to_sfixed(-0.9677,1,L_SIZE),
				to_sfixed(-0.9676,1,L_SIZE),
				to_sfixed(-0.9676,1,L_SIZE),
				to_sfixed(-0.9676,1,L_SIZE),
				to_sfixed(-0.9676,1,L_SIZE),
				to_sfixed(-0.9675,1,L_SIZE),
				to_sfixed(-0.9675,1,L_SIZE),
				to_sfixed(-0.9675,1,L_SIZE),
				to_sfixed(-0.9675,1,L_SIZE),
				to_sfixed(-0.9674,1,L_SIZE),
				to_sfixed(-0.9674,1,L_SIZE),
				to_sfixed(-0.9674,1,L_SIZE),
				to_sfixed(-0.9674,1,L_SIZE),
				to_sfixed(-0.9674,1,L_SIZE),
				to_sfixed(-0.9673,1,L_SIZE),
				to_sfixed(-0.9673,1,L_SIZE),
				to_sfixed(-0.9673,1,L_SIZE),
				to_sfixed(-0.9673,1,L_SIZE),
				to_sfixed(-0.9672,1,L_SIZE),
				to_sfixed(-0.9672,1,L_SIZE),
				to_sfixed(-0.9672,1,L_SIZE),
				to_sfixed(-0.9672,1,L_SIZE),
				to_sfixed(-0.9671,1,L_SIZE),
				to_sfixed(-0.9671,1,L_SIZE),
				to_sfixed(-0.9671,1,L_SIZE),
				to_sfixed(-0.9671,1,L_SIZE),
				to_sfixed(-0.9670,1,L_SIZE),
				to_sfixed(-0.9670,1,L_SIZE),
				to_sfixed(-0.9670,1,L_SIZE),
				to_sfixed(-0.9670,1,L_SIZE),
				to_sfixed(-0.9669,1,L_SIZE),
				to_sfixed(-0.9669,1,L_SIZE),
				to_sfixed(-0.9669,1,L_SIZE),
				to_sfixed(-0.9669,1,L_SIZE),
				to_sfixed(-0.9669,1,L_SIZE),
				to_sfixed(-0.9668,1,L_SIZE),
				to_sfixed(-0.9668,1,L_SIZE),
				to_sfixed(-0.9668,1,L_SIZE),
				to_sfixed(-0.9668,1,L_SIZE),
				to_sfixed(-0.9667,1,L_SIZE),
				to_sfixed(-0.9667,1,L_SIZE),
				to_sfixed(-0.9667,1,L_SIZE),
				to_sfixed(-0.9667,1,L_SIZE),
				to_sfixed(-0.9666,1,L_SIZE),
				to_sfixed(-0.9666,1,L_SIZE),
				to_sfixed(-0.9666,1,L_SIZE),
				to_sfixed(-0.9666,1,L_SIZE),
				to_sfixed(-0.9665,1,L_SIZE),
				to_sfixed(-0.9665,1,L_SIZE),
				to_sfixed(-0.9665,1,L_SIZE),
				to_sfixed(-0.9665,1,L_SIZE),
				to_sfixed(-0.9664,1,L_SIZE),
				to_sfixed(-0.9664,1,L_SIZE),
				to_sfixed(-0.9664,1,L_SIZE),
				to_sfixed(-0.9664,1,L_SIZE),
				to_sfixed(-0.9663,1,L_SIZE),
				to_sfixed(-0.9663,1,L_SIZE),
				to_sfixed(-0.9663,1,L_SIZE),
				to_sfixed(-0.9663,1,L_SIZE),
				to_sfixed(-0.9663,1,L_SIZE),
				to_sfixed(-0.9662,1,L_SIZE),
				to_sfixed(-0.9662,1,L_SIZE),
				to_sfixed(-0.9662,1,L_SIZE),
				to_sfixed(-0.9662,1,L_SIZE),
				to_sfixed(-0.9661,1,L_SIZE),
				to_sfixed(-0.9661,1,L_SIZE),
				to_sfixed(-0.9661,1,L_SIZE),
				to_sfixed(-0.9661,1,L_SIZE),
				to_sfixed(-0.9660,1,L_SIZE),
				to_sfixed(-0.9660,1,L_SIZE),
				to_sfixed(-0.9660,1,L_SIZE),
				to_sfixed(-0.9660,1,L_SIZE),
				to_sfixed(-0.9659,1,L_SIZE),
				to_sfixed(-0.9659,1,L_SIZE),
				to_sfixed(-0.9659,1,L_SIZE),
				to_sfixed(-0.9659,1,L_SIZE),
				to_sfixed(-0.9658,1,L_SIZE),
				to_sfixed(-0.9658,1,L_SIZE),
				to_sfixed(-0.9658,1,L_SIZE),
				to_sfixed(-0.9658,1,L_SIZE),
				to_sfixed(-0.9657,1,L_SIZE),
				to_sfixed(-0.9657,1,L_SIZE),
				to_sfixed(-0.9657,1,L_SIZE),
				to_sfixed(-0.9657,1,L_SIZE),
				to_sfixed(-0.9656,1,L_SIZE),
				to_sfixed(-0.9656,1,L_SIZE),
				to_sfixed(-0.9656,1,L_SIZE),
				to_sfixed(-0.9656,1,L_SIZE),
				to_sfixed(-0.9655,1,L_SIZE),
				to_sfixed(-0.9655,1,L_SIZE),
				to_sfixed(-0.9655,1,L_SIZE),
				to_sfixed(-0.9655,1,L_SIZE),
				to_sfixed(-0.9654,1,L_SIZE),
				to_sfixed(-0.9654,1,L_SIZE),
				to_sfixed(-0.9654,1,L_SIZE),
				to_sfixed(-0.9654,1,L_SIZE),
				to_sfixed(-0.9653,1,L_SIZE),
				to_sfixed(-0.9653,1,L_SIZE),
				to_sfixed(-0.9653,1,L_SIZE),
				to_sfixed(-0.9653,1,L_SIZE),
				to_sfixed(-0.9652,1,L_SIZE),
				to_sfixed(-0.9652,1,L_SIZE),
				to_sfixed(-0.9652,1,L_SIZE),
				to_sfixed(-0.9652,1,L_SIZE),
				to_sfixed(-0.9651,1,L_SIZE),
				to_sfixed(-0.9651,1,L_SIZE),
				to_sfixed(-0.9651,1,L_SIZE),
				to_sfixed(-0.9651,1,L_SIZE),
				to_sfixed(-0.9650,1,L_SIZE),
				to_sfixed(-0.9650,1,L_SIZE),
				to_sfixed(-0.9650,1,L_SIZE),
				to_sfixed(-0.9650,1,L_SIZE),
				to_sfixed(-0.9649,1,L_SIZE),
				to_sfixed(-0.9649,1,L_SIZE),
				to_sfixed(-0.9649,1,L_SIZE),
				to_sfixed(-0.9649,1,L_SIZE),
				to_sfixed(-0.9648,1,L_SIZE),
				to_sfixed(-0.9648,1,L_SIZE),
				to_sfixed(-0.9648,1,L_SIZE),
				to_sfixed(-0.9648,1,L_SIZE),
				to_sfixed(-0.9647,1,L_SIZE),
				to_sfixed(-0.9647,1,L_SIZE),
				to_sfixed(-0.9647,1,L_SIZE),
				to_sfixed(-0.9647,1,L_SIZE),
				to_sfixed(-0.9646,1,L_SIZE),
				to_sfixed(-0.9646,1,L_SIZE),
				to_sfixed(-0.9646,1,L_SIZE),
				to_sfixed(-0.9646,1,L_SIZE),
				to_sfixed(-0.9645,1,L_SIZE),
				to_sfixed(-0.9645,1,L_SIZE),
				to_sfixed(-0.9645,1,L_SIZE),
				to_sfixed(-0.9645,1,L_SIZE),
				to_sfixed(-0.9644,1,L_SIZE),
				to_sfixed(-0.9644,1,L_SIZE),
				to_sfixed(-0.9644,1,L_SIZE),
				to_sfixed(-0.9644,1,L_SIZE),
				to_sfixed(-0.9643,1,L_SIZE),
				to_sfixed(-0.9643,1,L_SIZE),
				to_sfixed(-0.9643,1,L_SIZE),
				to_sfixed(-0.9643,1,L_SIZE),
				to_sfixed(-0.9642,1,L_SIZE),
				to_sfixed(-0.9642,1,L_SIZE),
				to_sfixed(-0.9642,1,L_SIZE),
				to_sfixed(-0.9641,1,L_SIZE),
				to_sfixed(-0.9641,1,L_SIZE),
				to_sfixed(-0.9641,1,L_SIZE),
				to_sfixed(-0.9641,1,L_SIZE),
				to_sfixed(-0.9640,1,L_SIZE),
				to_sfixed(-0.9640,1,L_SIZE),
				to_sfixed(-0.9640,1,L_SIZE),
				to_sfixed(-0.9640,1,L_SIZE),
				to_sfixed(-0.9639,1,L_SIZE),
				to_sfixed(-0.9639,1,L_SIZE),
				to_sfixed(-0.9639,1,L_SIZE),
				to_sfixed(-0.9639,1,L_SIZE),
				to_sfixed(-0.9638,1,L_SIZE),
				to_sfixed(-0.9638,1,L_SIZE),
				to_sfixed(-0.9638,1,L_SIZE),
				to_sfixed(-0.9638,1,L_SIZE),
				to_sfixed(-0.9637,1,L_SIZE),
				to_sfixed(-0.9637,1,L_SIZE),
				to_sfixed(-0.9637,1,L_SIZE),
				to_sfixed(-0.9637,1,L_SIZE),
				to_sfixed(-0.9636,1,L_SIZE),
				to_sfixed(-0.9636,1,L_SIZE),
				to_sfixed(-0.9636,1,L_SIZE),
				to_sfixed(-0.9636,1,L_SIZE),
				to_sfixed(-0.9635,1,L_SIZE),
				to_sfixed(-0.9635,1,L_SIZE),
				to_sfixed(-0.9635,1,L_SIZE),
				to_sfixed(-0.9634,1,L_SIZE),
				to_sfixed(-0.9634,1,L_SIZE),
				to_sfixed(-0.9634,1,L_SIZE),
				to_sfixed(-0.9634,1,L_SIZE),
				to_sfixed(-0.9633,1,L_SIZE),
				to_sfixed(-0.9633,1,L_SIZE),
				to_sfixed(-0.9633,1,L_SIZE),
				to_sfixed(-0.9633,1,L_SIZE),
				to_sfixed(-0.9632,1,L_SIZE),
				to_sfixed(-0.9632,1,L_SIZE),
				to_sfixed(-0.9632,1,L_SIZE),
				to_sfixed(-0.9632,1,L_SIZE),
				to_sfixed(-0.9631,1,L_SIZE),
				to_sfixed(-0.9631,1,L_SIZE),
				to_sfixed(-0.9631,1,L_SIZE),
				to_sfixed(-0.9630,1,L_SIZE),
				to_sfixed(-0.9630,1,L_SIZE),
				to_sfixed(-0.9630,1,L_SIZE),
				to_sfixed(-0.9630,1,L_SIZE),
				to_sfixed(-0.9629,1,L_SIZE),
				to_sfixed(-0.9629,1,L_SIZE),
				to_sfixed(-0.9629,1,L_SIZE),
				to_sfixed(-0.9629,1,L_SIZE),
				to_sfixed(-0.9628,1,L_SIZE),
				to_sfixed(-0.9628,1,L_SIZE),
				to_sfixed(-0.9628,1,L_SIZE),
				to_sfixed(-0.9628,1,L_SIZE),
				to_sfixed(-0.9627,1,L_SIZE),
				to_sfixed(-0.9627,1,L_SIZE),
				to_sfixed(-0.9627,1,L_SIZE),
				to_sfixed(-0.9626,1,L_SIZE),
				to_sfixed(-0.9626,1,L_SIZE),
				to_sfixed(-0.9626,1,L_SIZE),
				to_sfixed(-0.9626,1,L_SIZE),
				to_sfixed(-0.9625,1,L_SIZE),
				to_sfixed(-0.9625,1,L_SIZE),
				to_sfixed(-0.9625,1,L_SIZE),
				to_sfixed(-0.9625,1,L_SIZE),
				to_sfixed(-0.9624,1,L_SIZE),
				to_sfixed(-0.9624,1,L_SIZE),
				to_sfixed(-0.9624,1,L_SIZE),
				to_sfixed(-0.9624,1,L_SIZE),
				to_sfixed(-0.9623,1,L_SIZE),
				to_sfixed(-0.9623,1,L_SIZE),
				to_sfixed(-0.9623,1,L_SIZE),
				to_sfixed(-0.9622,1,L_SIZE),
				to_sfixed(-0.9622,1,L_SIZE),
				to_sfixed(-0.9622,1,L_SIZE),
				to_sfixed(-0.9622,1,L_SIZE),
				to_sfixed(-0.9621,1,L_SIZE),
				to_sfixed(-0.9621,1,L_SIZE),
				to_sfixed(-0.9621,1,L_SIZE),
				to_sfixed(-0.9621,1,L_SIZE),
				to_sfixed(-0.9620,1,L_SIZE),
				to_sfixed(-0.9620,1,L_SIZE),
				to_sfixed(-0.9620,1,L_SIZE),
				to_sfixed(-0.9619,1,L_SIZE),
				to_sfixed(-0.9619,1,L_SIZE),
				to_sfixed(-0.9619,1,L_SIZE),
				to_sfixed(-0.9619,1,L_SIZE),
				to_sfixed(-0.9618,1,L_SIZE),
				to_sfixed(-0.9618,1,L_SIZE),
				to_sfixed(-0.9618,1,L_SIZE),
				to_sfixed(-0.9618,1,L_SIZE),
				to_sfixed(-0.9617,1,L_SIZE),
				to_sfixed(-0.9617,1,L_SIZE),
				to_sfixed(-0.9617,1,L_SIZE),
				to_sfixed(-0.9616,1,L_SIZE),
				to_sfixed(-0.9616,1,L_SIZE),
				to_sfixed(-0.9616,1,L_SIZE),
				to_sfixed(-0.9616,1,L_SIZE),
				to_sfixed(-0.9615,1,L_SIZE),
				to_sfixed(-0.9615,1,L_SIZE),
				to_sfixed(-0.9615,1,L_SIZE),
				to_sfixed(-0.9614,1,L_SIZE),
				to_sfixed(-0.9614,1,L_SIZE),
				to_sfixed(-0.9614,1,L_SIZE),
				to_sfixed(-0.9614,1,L_SIZE),
				to_sfixed(-0.9613,1,L_SIZE),
				to_sfixed(-0.9613,1,L_SIZE),
				to_sfixed(-0.9613,1,L_SIZE),
				to_sfixed(-0.9613,1,L_SIZE),
				to_sfixed(-0.9612,1,L_SIZE),
				to_sfixed(-0.9612,1,L_SIZE),
				to_sfixed(-0.9612,1,L_SIZE),
				to_sfixed(-0.9611,1,L_SIZE),
				to_sfixed(-0.9611,1,L_SIZE),
				to_sfixed(-0.9611,1,L_SIZE),
				to_sfixed(-0.9611,1,L_SIZE),
				to_sfixed(-0.9610,1,L_SIZE),
				to_sfixed(-0.9610,1,L_SIZE),
				to_sfixed(-0.9610,1,L_SIZE),
				to_sfixed(-0.9609,1,L_SIZE),
				to_sfixed(-0.9609,1,L_SIZE),
				to_sfixed(-0.9609,1,L_SIZE),
				to_sfixed(-0.9609,1,L_SIZE),
				to_sfixed(-0.9608,1,L_SIZE),
				to_sfixed(-0.9608,1,L_SIZE),
				to_sfixed(-0.9608,1,L_SIZE),
				to_sfixed(-0.9608,1,L_SIZE),
				to_sfixed(-0.9607,1,L_SIZE),
				to_sfixed(-0.9607,1,L_SIZE),
				to_sfixed(-0.9607,1,L_SIZE),
				to_sfixed(-0.9606,1,L_SIZE),
				to_sfixed(-0.9606,1,L_SIZE),
				to_sfixed(-0.9606,1,L_SIZE),
				to_sfixed(-0.9606,1,L_SIZE),
				to_sfixed(-0.9605,1,L_SIZE),
				to_sfixed(-0.9605,1,L_SIZE),
				to_sfixed(-0.9605,1,L_SIZE),
				to_sfixed(-0.9604,1,L_SIZE),
				to_sfixed(-0.9604,1,L_SIZE),
				to_sfixed(-0.9604,1,L_SIZE),
				to_sfixed(-0.9604,1,L_SIZE),
				to_sfixed(-0.9603,1,L_SIZE),
				to_sfixed(-0.9603,1,L_SIZE),
				to_sfixed(-0.9603,1,L_SIZE),
				to_sfixed(-0.9602,1,L_SIZE),
				to_sfixed(-0.9602,1,L_SIZE),
				to_sfixed(-0.9602,1,L_SIZE),
				to_sfixed(-0.9602,1,L_SIZE),
				to_sfixed(-0.9601,1,L_SIZE),
				to_sfixed(-0.9601,1,L_SIZE),
				to_sfixed(-0.9601,1,L_SIZE),
				to_sfixed(-0.9600,1,L_SIZE),
				to_sfixed(-0.9600,1,L_SIZE),
				to_sfixed(-0.9600,1,L_SIZE),
				to_sfixed(-0.9600,1,L_SIZE),
				to_sfixed(-0.9599,1,L_SIZE),
				to_sfixed(-0.9599,1,L_SIZE),
				to_sfixed(-0.9599,1,L_SIZE),
				to_sfixed(-0.9598,1,L_SIZE),
				to_sfixed(-0.9598,1,L_SIZE),
				to_sfixed(-0.9598,1,L_SIZE),
				to_sfixed(-0.9598,1,L_SIZE),
				to_sfixed(-0.9597,1,L_SIZE),
				to_sfixed(-0.9597,1,L_SIZE),
				to_sfixed(-0.9597,1,L_SIZE),
				to_sfixed(-0.9596,1,L_SIZE),
				to_sfixed(-0.9596,1,L_SIZE),
				to_sfixed(-0.9596,1,L_SIZE),
				to_sfixed(-0.9595,1,L_SIZE),
				to_sfixed(-0.9595,1,L_SIZE),
				to_sfixed(-0.9595,1,L_SIZE),
				to_sfixed(-0.9595,1,L_SIZE),
				to_sfixed(-0.9594,1,L_SIZE),
				to_sfixed(-0.9594,1,L_SIZE),
				to_sfixed(-0.9594,1,L_SIZE),
				to_sfixed(-0.9593,1,L_SIZE),
				to_sfixed(-0.9593,1,L_SIZE),
				to_sfixed(-0.9593,1,L_SIZE),
				to_sfixed(-0.9593,1,L_SIZE),
				to_sfixed(-0.9592,1,L_SIZE),
				to_sfixed(-0.9592,1,L_SIZE),
				to_sfixed(-0.9592,1,L_SIZE),
				to_sfixed(-0.9591,1,L_SIZE),
				to_sfixed(-0.9591,1,L_SIZE),
				to_sfixed(-0.9591,1,L_SIZE),
				to_sfixed(-0.9591,1,L_SIZE),
				to_sfixed(-0.9590,1,L_SIZE),
				to_sfixed(-0.9590,1,L_SIZE),
				to_sfixed(-0.9590,1,L_SIZE),
				to_sfixed(-0.9589,1,L_SIZE),
				to_sfixed(-0.9589,1,L_SIZE),
				to_sfixed(-0.9589,1,L_SIZE),
				to_sfixed(-0.9588,1,L_SIZE),
				to_sfixed(-0.9588,1,L_SIZE),
				to_sfixed(-0.9588,1,L_SIZE),
				to_sfixed(-0.9588,1,L_SIZE),
				to_sfixed(-0.9587,1,L_SIZE),
				to_sfixed(-0.9587,1,L_SIZE),
				to_sfixed(-0.9587,1,L_SIZE),
				to_sfixed(-0.9586,1,L_SIZE),
				to_sfixed(-0.9586,1,L_SIZE),
				to_sfixed(-0.9586,1,L_SIZE),
				to_sfixed(-0.9585,1,L_SIZE),
				to_sfixed(-0.9585,1,L_SIZE),
				to_sfixed(-0.9585,1,L_SIZE),
				to_sfixed(-0.9585,1,L_SIZE),
				to_sfixed(-0.9584,1,L_SIZE),
				to_sfixed(-0.9584,1,L_SIZE),
				to_sfixed(-0.9584,1,L_SIZE),
				to_sfixed(-0.9583,1,L_SIZE),
				to_sfixed(-0.9583,1,L_SIZE),
				to_sfixed(-0.9583,1,L_SIZE),
				to_sfixed(-0.9583,1,L_SIZE),
				to_sfixed(-0.9582,1,L_SIZE),
				to_sfixed(-0.9582,1,L_SIZE),
				to_sfixed(-0.9582,1,L_SIZE),
				to_sfixed(-0.9581,1,L_SIZE),
				to_sfixed(-0.9581,1,L_SIZE),
				to_sfixed(-0.9581,1,L_SIZE),
				to_sfixed(-0.9580,1,L_SIZE),
				to_sfixed(-0.9580,1,L_SIZE),
				to_sfixed(-0.9580,1,L_SIZE),
				to_sfixed(-0.9580,1,L_SIZE),
				to_sfixed(-0.9579,1,L_SIZE),
				to_sfixed(-0.9579,1,L_SIZE),
				to_sfixed(-0.9579,1,L_SIZE),
				to_sfixed(-0.9578,1,L_SIZE),
				to_sfixed(-0.9578,1,L_SIZE),
				to_sfixed(-0.9578,1,L_SIZE),
				to_sfixed(-0.9577,1,L_SIZE),
				to_sfixed(-0.9577,1,L_SIZE),
				to_sfixed(-0.9577,1,L_SIZE),
				to_sfixed(-0.9576,1,L_SIZE),
				to_sfixed(-0.9576,1,L_SIZE),
				to_sfixed(-0.9576,1,L_SIZE),
				to_sfixed(-0.9576,1,L_SIZE),
				to_sfixed(-0.9575,1,L_SIZE),
				to_sfixed(-0.9575,1,L_SIZE),
				to_sfixed(-0.9575,1,L_SIZE),
				to_sfixed(-0.9574,1,L_SIZE),
				to_sfixed(-0.9574,1,L_SIZE),
				to_sfixed(-0.9574,1,L_SIZE),
				to_sfixed(-0.9573,1,L_SIZE),
				to_sfixed(-0.9573,1,L_SIZE),
				to_sfixed(-0.9573,1,L_SIZE),
				to_sfixed(-0.9573,1,L_SIZE),
				to_sfixed(-0.9572,1,L_SIZE),
				to_sfixed(-0.9572,1,L_SIZE),
				to_sfixed(-0.9572,1,L_SIZE),
				to_sfixed(-0.9571,1,L_SIZE),
				to_sfixed(-0.9571,1,L_SIZE),
				to_sfixed(-0.9571,1,L_SIZE),
				to_sfixed(-0.9570,1,L_SIZE),
				to_sfixed(-0.9570,1,L_SIZE),
				to_sfixed(-0.9570,1,L_SIZE),
				to_sfixed(-0.9569,1,L_SIZE),
				to_sfixed(-0.9569,1,L_SIZE),
				to_sfixed(-0.9569,1,L_SIZE),
				to_sfixed(-0.9569,1,L_SIZE),
				to_sfixed(-0.9568,1,L_SIZE),
				to_sfixed(-0.9568,1,L_SIZE),
				to_sfixed(-0.9568,1,L_SIZE),
				to_sfixed(-0.9567,1,L_SIZE),
				to_sfixed(-0.9567,1,L_SIZE),
				to_sfixed(-0.9567,1,L_SIZE),
				to_sfixed(-0.9566,1,L_SIZE),
				to_sfixed(-0.9566,1,L_SIZE),
				to_sfixed(-0.9566,1,L_SIZE),
				to_sfixed(-0.9565,1,L_SIZE),
				to_sfixed(-0.9565,1,L_SIZE),
				to_sfixed(-0.9565,1,L_SIZE),
				to_sfixed(-0.9564,1,L_SIZE),
				to_sfixed(-0.9564,1,L_SIZE),
				to_sfixed(-0.9564,1,L_SIZE),
				to_sfixed(-0.9564,1,L_SIZE),
				to_sfixed(-0.9563,1,L_SIZE),
				to_sfixed(-0.9563,1,L_SIZE),
				to_sfixed(-0.9563,1,L_SIZE),
				to_sfixed(-0.9562,1,L_SIZE),
				to_sfixed(-0.9562,1,L_SIZE),
				to_sfixed(-0.9562,1,L_SIZE),
				to_sfixed(-0.9561,1,L_SIZE),
				to_sfixed(-0.9561,1,L_SIZE),
				to_sfixed(-0.9561,1,L_SIZE),
				to_sfixed(-0.9560,1,L_SIZE),
				to_sfixed(-0.9560,1,L_SIZE),
				to_sfixed(-0.9560,1,L_SIZE),
				to_sfixed(-0.9559,1,L_SIZE),
				to_sfixed(-0.9559,1,L_SIZE),
				to_sfixed(-0.9559,1,L_SIZE),
				to_sfixed(-0.9559,1,L_SIZE),
				to_sfixed(-0.9558,1,L_SIZE),
				to_sfixed(-0.9558,1,L_SIZE),
				to_sfixed(-0.9558,1,L_SIZE),
				to_sfixed(-0.9557,1,L_SIZE),
				to_sfixed(-0.9557,1,L_SIZE),
				to_sfixed(-0.9557,1,L_SIZE),
				to_sfixed(-0.9556,1,L_SIZE),
				to_sfixed(-0.9556,1,L_SIZE),
				to_sfixed(-0.9556,1,L_SIZE),
				to_sfixed(-0.9555,1,L_SIZE),
				to_sfixed(-0.9555,1,L_SIZE),
				to_sfixed(-0.9555,1,L_SIZE),
				to_sfixed(-0.9554,1,L_SIZE),
				to_sfixed(-0.9554,1,L_SIZE),
				to_sfixed(-0.9554,1,L_SIZE),
				to_sfixed(-0.9553,1,L_SIZE),
				to_sfixed(-0.9553,1,L_SIZE),
				to_sfixed(-0.9553,1,L_SIZE),
				to_sfixed(-0.9552,1,L_SIZE),
				to_sfixed(-0.9552,1,L_SIZE),
				to_sfixed(-0.9552,1,L_SIZE),
				to_sfixed(-0.9552,1,L_SIZE),
				to_sfixed(-0.9551,1,L_SIZE),
				to_sfixed(-0.9551,1,L_SIZE),
				to_sfixed(-0.9551,1,L_SIZE),
				to_sfixed(-0.9550,1,L_SIZE),
				to_sfixed(-0.9550,1,L_SIZE),
				to_sfixed(-0.9550,1,L_SIZE),
				to_sfixed(-0.9549,1,L_SIZE),
				to_sfixed(-0.9549,1,L_SIZE),
				to_sfixed(-0.9549,1,L_SIZE),
				to_sfixed(-0.9548,1,L_SIZE),
				to_sfixed(-0.9548,1,L_SIZE),
				to_sfixed(-0.9548,1,L_SIZE),
				to_sfixed(-0.9547,1,L_SIZE),
				to_sfixed(-0.9547,1,L_SIZE),
				to_sfixed(-0.9547,1,L_SIZE),
				to_sfixed(-0.9546,1,L_SIZE),
				to_sfixed(-0.9546,1,L_SIZE),
				to_sfixed(-0.9546,1,L_SIZE),
				to_sfixed(-0.9545,1,L_SIZE),
				to_sfixed(-0.9545,1,L_SIZE),
				to_sfixed(-0.9545,1,L_SIZE),
				to_sfixed(-0.9544,1,L_SIZE),
				to_sfixed(-0.9544,1,L_SIZE),
				to_sfixed(-0.9544,1,L_SIZE),
				to_sfixed(-0.9543,1,L_SIZE),
				to_sfixed(-0.9543,1,L_SIZE),
				to_sfixed(-0.9543,1,L_SIZE),
				to_sfixed(-0.9542,1,L_SIZE),
				to_sfixed(-0.9542,1,L_SIZE),
				to_sfixed(-0.9542,1,L_SIZE),
				to_sfixed(-0.9541,1,L_SIZE),
				to_sfixed(-0.9541,1,L_SIZE),
				to_sfixed(-0.9541,1,L_SIZE),
				to_sfixed(-0.9540,1,L_SIZE),
				to_sfixed(-0.9540,1,L_SIZE),
				to_sfixed(-0.9540,1,L_SIZE),
				to_sfixed(-0.9539,1,L_SIZE),
				to_sfixed(-0.9539,1,L_SIZE),
				to_sfixed(-0.9539,1,L_SIZE),
				to_sfixed(-0.9538,1,L_SIZE),
				to_sfixed(-0.9538,1,L_SIZE),
				to_sfixed(-0.9538,1,L_SIZE),
				to_sfixed(-0.9537,1,L_SIZE),
				to_sfixed(-0.9537,1,L_SIZE),
				to_sfixed(-0.9537,1,L_SIZE),
				to_sfixed(-0.9536,1,L_SIZE),
				to_sfixed(-0.9536,1,L_SIZE),
				to_sfixed(-0.9536,1,L_SIZE),
				to_sfixed(-0.9535,1,L_SIZE),
				to_sfixed(-0.9535,1,L_SIZE),
				to_sfixed(-0.9535,1,L_SIZE),
				to_sfixed(-0.9534,1,L_SIZE),
				to_sfixed(-0.9534,1,L_SIZE),
				to_sfixed(-0.9534,1,L_SIZE),
				to_sfixed(-0.9533,1,L_SIZE),
				to_sfixed(-0.9533,1,L_SIZE),
				to_sfixed(-0.9533,1,L_SIZE),
				to_sfixed(-0.9532,1,L_SIZE),
				to_sfixed(-0.9532,1,L_SIZE),
				to_sfixed(-0.9532,1,L_SIZE),
				to_sfixed(-0.9531,1,L_SIZE),
				to_sfixed(-0.9531,1,L_SIZE),
				to_sfixed(-0.9531,1,L_SIZE),
				to_sfixed(-0.9530,1,L_SIZE),
				to_sfixed(-0.9530,1,L_SIZE),
				to_sfixed(-0.9530,1,L_SIZE),
				to_sfixed(-0.9529,1,L_SIZE),
				to_sfixed(-0.9529,1,L_SIZE),
				to_sfixed(-0.9529,1,L_SIZE),
				to_sfixed(-0.9528,1,L_SIZE),
				to_sfixed(-0.9528,1,L_SIZE),
				to_sfixed(-0.9528,1,L_SIZE),
				to_sfixed(-0.9527,1,L_SIZE),
				to_sfixed(-0.9527,1,L_SIZE),
				to_sfixed(-0.9527,1,L_SIZE),
				to_sfixed(-0.9526,1,L_SIZE),
				to_sfixed(-0.9526,1,L_SIZE),
				to_sfixed(-0.9526,1,L_SIZE),
				to_sfixed(-0.9525,1,L_SIZE),
				to_sfixed(-0.9525,1,L_SIZE),
				to_sfixed(-0.9525,1,L_SIZE),
				to_sfixed(-0.9524,1,L_SIZE),
				to_sfixed(-0.9524,1,L_SIZE),
				to_sfixed(-0.9524,1,L_SIZE),
				to_sfixed(-0.9523,1,L_SIZE),
				to_sfixed(-0.9523,1,L_SIZE),
				to_sfixed(-0.9523,1,L_SIZE),
				to_sfixed(-0.9522,1,L_SIZE),
				to_sfixed(-0.9522,1,L_SIZE),
				to_sfixed(-0.9522,1,L_SIZE),
				to_sfixed(-0.9521,1,L_SIZE),
				to_sfixed(-0.9521,1,L_SIZE),
				to_sfixed(-0.9521,1,L_SIZE),
				to_sfixed(-0.9520,1,L_SIZE),
				to_sfixed(-0.9520,1,L_SIZE),
				to_sfixed(-0.9520,1,L_SIZE),
				to_sfixed(-0.9519,1,L_SIZE),
				to_sfixed(-0.9519,1,L_SIZE),
				to_sfixed(-0.9519,1,L_SIZE),
				to_sfixed(-0.9518,1,L_SIZE),
				to_sfixed(-0.9518,1,L_SIZE),
				to_sfixed(-0.9518,1,L_SIZE),
				to_sfixed(-0.9517,1,L_SIZE),
				to_sfixed(-0.9517,1,L_SIZE),
				to_sfixed(-0.9517,1,L_SIZE),
				to_sfixed(-0.9516,1,L_SIZE),
				to_sfixed(-0.9516,1,L_SIZE),
				to_sfixed(-0.9515,1,L_SIZE),
				to_sfixed(-0.9515,1,L_SIZE),
				to_sfixed(-0.9515,1,L_SIZE),
				to_sfixed(-0.9514,1,L_SIZE),
				to_sfixed(-0.9514,1,L_SIZE),
				to_sfixed(-0.9514,1,L_SIZE),
				to_sfixed(-0.9513,1,L_SIZE),
				to_sfixed(-0.9513,1,L_SIZE),
				to_sfixed(-0.9513,1,L_SIZE),
				to_sfixed(-0.9512,1,L_SIZE),
				to_sfixed(-0.9512,1,L_SIZE),
				to_sfixed(-0.9512,1,L_SIZE),
				to_sfixed(-0.9511,1,L_SIZE),
				to_sfixed(-0.9511,1,L_SIZE),
				to_sfixed(-0.9511,1,L_SIZE),
				to_sfixed(-0.9510,1,L_SIZE),
				to_sfixed(-0.9510,1,L_SIZE),
				to_sfixed(-0.9510,1,L_SIZE),
				to_sfixed(-0.9509,1,L_SIZE),
				to_sfixed(-0.9509,1,L_SIZE),
				to_sfixed(-0.9509,1,L_SIZE),
				to_sfixed(-0.9508,1,L_SIZE),
				to_sfixed(-0.9508,1,L_SIZE),
				to_sfixed(-0.9507,1,L_SIZE),
				to_sfixed(-0.9507,1,L_SIZE),
				to_sfixed(-0.9507,1,L_SIZE),
				to_sfixed(-0.9506,1,L_SIZE),
				to_sfixed(-0.9506,1,L_SIZE),
				to_sfixed(-0.9506,1,L_SIZE),
				to_sfixed(-0.9505,1,L_SIZE),
				to_sfixed(-0.9505,1,L_SIZE),
				to_sfixed(-0.9505,1,L_SIZE),
				to_sfixed(-0.9504,1,L_SIZE),
				to_sfixed(-0.9504,1,L_SIZE),
				to_sfixed(-0.9504,1,L_SIZE),
				to_sfixed(-0.9503,1,L_SIZE),
				to_sfixed(-0.9503,1,L_SIZE),
				to_sfixed(-0.9502,1,L_SIZE),
				to_sfixed(-0.9502,1,L_SIZE),
				to_sfixed(-0.9502,1,L_SIZE),
				to_sfixed(-0.9501,1,L_SIZE),
				to_sfixed(-0.9501,1,L_SIZE),
				to_sfixed(-0.9501,1,L_SIZE),
				to_sfixed(-0.9500,1,L_SIZE),
				to_sfixed(-0.9500,1,L_SIZE),
				to_sfixed(-0.9500,1,L_SIZE),
				to_sfixed(-0.9499,1,L_SIZE),
				to_sfixed(-0.9499,1,L_SIZE),
				to_sfixed(-0.9499,1,L_SIZE),
				to_sfixed(-0.9498,1,L_SIZE),
				to_sfixed(-0.9498,1,L_SIZE),
				to_sfixed(-0.9498,1,L_SIZE),
				to_sfixed(-0.9497,1,L_SIZE),
				to_sfixed(-0.9497,1,L_SIZE),
				to_sfixed(-0.9496,1,L_SIZE),
				to_sfixed(-0.9496,1,L_SIZE),
				to_sfixed(-0.9496,1,L_SIZE),
				to_sfixed(-0.9495,1,L_SIZE),
				to_sfixed(-0.9495,1,L_SIZE),
				to_sfixed(-0.9495,1,L_SIZE),
				to_sfixed(-0.9494,1,L_SIZE),
				to_sfixed(-0.9494,1,L_SIZE),
				to_sfixed(-0.9494,1,L_SIZE),
				to_sfixed(-0.9493,1,L_SIZE),
				to_sfixed(-0.9493,1,L_SIZE),
				to_sfixed(-0.9492,1,L_SIZE),
				to_sfixed(-0.9492,1,L_SIZE),
				to_sfixed(-0.9492,1,L_SIZE),
				to_sfixed(-0.9491,1,L_SIZE),
				to_sfixed(-0.9491,1,L_SIZE),
				to_sfixed(-0.9491,1,L_SIZE),
				to_sfixed(-0.9490,1,L_SIZE),
				to_sfixed(-0.9490,1,L_SIZE),
				to_sfixed(-0.9490,1,L_SIZE),
				to_sfixed(-0.9489,1,L_SIZE),
				to_sfixed(-0.9489,1,L_SIZE),
				to_sfixed(-0.9488,1,L_SIZE),
				to_sfixed(-0.9488,1,L_SIZE),
				to_sfixed(-0.9488,1,L_SIZE),
				to_sfixed(-0.9487,1,L_SIZE),
				to_sfixed(-0.9487,1,L_SIZE),
				to_sfixed(-0.9487,1,L_SIZE),
				to_sfixed(-0.9486,1,L_SIZE),
				to_sfixed(-0.9486,1,L_SIZE),
				to_sfixed(-0.9486,1,L_SIZE),
				to_sfixed(-0.9485,1,L_SIZE),
				to_sfixed(-0.9485,1,L_SIZE),
				to_sfixed(-0.9484,1,L_SIZE),
				to_sfixed(-0.9484,1,L_SIZE),
				to_sfixed(-0.9484,1,L_SIZE),
				to_sfixed(-0.9483,1,L_SIZE),
				to_sfixed(-0.9483,1,L_SIZE),
				to_sfixed(-0.9483,1,L_SIZE),
				to_sfixed(-0.9482,1,L_SIZE),
				to_sfixed(-0.9482,1,L_SIZE),
				to_sfixed(-0.9481,1,L_SIZE),
				to_sfixed(-0.9481,1,L_SIZE),
				to_sfixed(-0.9481,1,L_SIZE),
				to_sfixed(-0.9480,1,L_SIZE),
				to_sfixed(-0.9480,1,L_SIZE),
				to_sfixed(-0.9480,1,L_SIZE),
				to_sfixed(-0.9479,1,L_SIZE),
				to_sfixed(-0.9479,1,L_SIZE),
				to_sfixed(-0.9479,1,L_SIZE),
				to_sfixed(-0.9478,1,L_SIZE),
				to_sfixed(-0.9478,1,L_SIZE),
				to_sfixed(-0.9477,1,L_SIZE),
				to_sfixed(-0.9477,1,L_SIZE),
				to_sfixed(-0.9477,1,L_SIZE),
				to_sfixed(-0.9476,1,L_SIZE),
				to_sfixed(-0.9476,1,L_SIZE),
				to_sfixed(-0.9476,1,L_SIZE),
				to_sfixed(-0.9475,1,L_SIZE),
				to_sfixed(-0.9475,1,L_SIZE),
				to_sfixed(-0.9474,1,L_SIZE),
				to_sfixed(-0.9474,1,L_SIZE),
				to_sfixed(-0.9474,1,L_SIZE),
				to_sfixed(-0.9473,1,L_SIZE),
				to_sfixed(-0.9473,1,L_SIZE),
				to_sfixed(-0.9473,1,L_SIZE),
				to_sfixed(-0.9472,1,L_SIZE),
				to_sfixed(-0.9472,1,L_SIZE),
				to_sfixed(-0.9471,1,L_SIZE),
				to_sfixed(-0.9471,1,L_SIZE),
				to_sfixed(-0.9471,1,L_SIZE),
				to_sfixed(-0.9470,1,L_SIZE),
				to_sfixed(-0.9470,1,L_SIZE),
				to_sfixed(-0.9469,1,L_SIZE),
				to_sfixed(-0.9469,1,L_SIZE),
				to_sfixed(-0.9469,1,L_SIZE),
				to_sfixed(-0.9468,1,L_SIZE),
				to_sfixed(-0.9468,1,L_SIZE),
				to_sfixed(-0.9468,1,L_SIZE),
				to_sfixed(-0.9467,1,L_SIZE),
				to_sfixed(-0.9467,1,L_SIZE),
				to_sfixed(-0.9466,1,L_SIZE),
				to_sfixed(-0.9466,1,L_SIZE),
				to_sfixed(-0.9466,1,L_SIZE),
				to_sfixed(-0.9465,1,L_SIZE),
				to_sfixed(-0.9465,1,L_SIZE),
				to_sfixed(-0.9465,1,L_SIZE),
				to_sfixed(-0.9464,1,L_SIZE),
				to_sfixed(-0.9464,1,L_SIZE),
				to_sfixed(-0.9463,1,L_SIZE),
				to_sfixed(-0.9463,1,L_SIZE),
				to_sfixed(-0.9463,1,L_SIZE),
				to_sfixed(-0.9462,1,L_SIZE),
				to_sfixed(-0.9462,1,L_SIZE),
				to_sfixed(-0.9461,1,L_SIZE),
				to_sfixed(-0.9461,1,L_SIZE),
				to_sfixed(-0.9461,1,L_SIZE),
				to_sfixed(-0.9460,1,L_SIZE),
				to_sfixed(-0.9460,1,L_SIZE),
				to_sfixed(-0.9460,1,L_SIZE),
				to_sfixed(-0.9459,1,L_SIZE),
				to_sfixed(-0.9459,1,L_SIZE),
				to_sfixed(-0.9458,1,L_SIZE),
				to_sfixed(-0.9458,1,L_SIZE),
				to_sfixed(-0.9458,1,L_SIZE),
				to_sfixed(-0.9457,1,L_SIZE),
				to_sfixed(-0.9457,1,L_SIZE),
				to_sfixed(-0.9456,1,L_SIZE),
				to_sfixed(-0.9456,1,L_SIZE),
				to_sfixed(-0.9456,1,L_SIZE),
				to_sfixed(-0.9455,1,L_SIZE),
				to_sfixed(-0.9455,1,L_SIZE),
				to_sfixed(-0.9455,1,L_SIZE),
				to_sfixed(-0.9454,1,L_SIZE),
				to_sfixed(-0.9454,1,L_SIZE),
				to_sfixed(-0.9453,1,L_SIZE),
				to_sfixed(-0.9453,1,L_SIZE),
				to_sfixed(-0.9453,1,L_SIZE),
				to_sfixed(-0.9452,1,L_SIZE),
				to_sfixed(-0.9452,1,L_SIZE),
				to_sfixed(-0.9451,1,L_SIZE),
				to_sfixed(-0.9451,1,L_SIZE),
				to_sfixed(-0.9451,1,L_SIZE),
				to_sfixed(-0.9450,1,L_SIZE),
				to_sfixed(-0.9450,1,L_SIZE),
				to_sfixed(-0.9449,1,L_SIZE),
				to_sfixed(-0.9449,1,L_SIZE),
				to_sfixed(-0.9449,1,L_SIZE),
				to_sfixed(-0.9448,1,L_SIZE),
				to_sfixed(-0.9448,1,L_SIZE),
				to_sfixed(-0.9448,1,L_SIZE),
				to_sfixed(-0.9447,1,L_SIZE),
				to_sfixed(-0.9447,1,L_SIZE),
				to_sfixed(-0.9446,1,L_SIZE),
				to_sfixed(-0.9446,1,L_SIZE),
				to_sfixed(-0.9446,1,L_SIZE),
				to_sfixed(-0.9445,1,L_SIZE),
				to_sfixed(-0.9445,1,L_SIZE),
				to_sfixed(-0.9444,1,L_SIZE),
				to_sfixed(-0.9444,1,L_SIZE),
				to_sfixed(-0.9444,1,L_SIZE),
				to_sfixed(-0.9443,1,L_SIZE),
				to_sfixed(-0.9443,1,L_SIZE),
				to_sfixed(-0.9442,1,L_SIZE),
				to_sfixed(-0.9442,1,L_SIZE),
				to_sfixed(-0.9442,1,L_SIZE),
				to_sfixed(-0.9441,1,L_SIZE),
				to_sfixed(-0.9441,1,L_SIZE),
				to_sfixed(-0.9440,1,L_SIZE),
				to_sfixed(-0.9440,1,L_SIZE),
				to_sfixed(-0.9440,1,L_SIZE),
				to_sfixed(-0.9439,1,L_SIZE),
				to_sfixed(-0.9439,1,L_SIZE),
				to_sfixed(-0.9438,1,L_SIZE),
				to_sfixed(-0.9438,1,L_SIZE),
				to_sfixed(-0.9438,1,L_SIZE),
				to_sfixed(-0.9437,1,L_SIZE),
				to_sfixed(-0.9437,1,L_SIZE),
				to_sfixed(-0.9436,1,L_SIZE),
				to_sfixed(-0.9436,1,L_SIZE),
				to_sfixed(-0.9436,1,L_SIZE),
				to_sfixed(-0.9435,1,L_SIZE),
				to_sfixed(-0.9435,1,L_SIZE),
				to_sfixed(-0.9434,1,L_SIZE),
				to_sfixed(-0.9434,1,L_SIZE),
				to_sfixed(-0.9434,1,L_SIZE),
				to_sfixed(-0.9433,1,L_SIZE),
				to_sfixed(-0.9433,1,L_SIZE),
				to_sfixed(-0.9432,1,L_SIZE),
				to_sfixed(-0.9432,1,L_SIZE),
				to_sfixed(-0.9432,1,L_SIZE),
				to_sfixed(-0.9431,1,L_SIZE),
				to_sfixed(-0.9431,1,L_SIZE),
				to_sfixed(-0.9430,1,L_SIZE),
				to_sfixed(-0.9430,1,L_SIZE),
				to_sfixed(-0.9430,1,L_SIZE),
				to_sfixed(-0.9429,1,L_SIZE),
				to_sfixed(-0.9429,1,L_SIZE),
				to_sfixed(-0.9428,1,L_SIZE),
				to_sfixed(-0.9428,1,L_SIZE),
				to_sfixed(-0.9427,1,L_SIZE),
				to_sfixed(-0.9427,1,L_SIZE),
				to_sfixed(-0.9427,1,L_SIZE),
				to_sfixed(-0.9426,1,L_SIZE),
				to_sfixed(-0.9426,1,L_SIZE),
				to_sfixed(-0.9425,1,L_SIZE),
				to_sfixed(-0.9425,1,L_SIZE),
				to_sfixed(-0.9425,1,L_SIZE),
				to_sfixed(-0.9424,1,L_SIZE),
				to_sfixed(-0.9424,1,L_SIZE),
				to_sfixed(-0.9423,1,L_SIZE),
				to_sfixed(-0.9423,1,L_SIZE),
				to_sfixed(-0.9423,1,L_SIZE),
				to_sfixed(-0.9422,1,L_SIZE),
				to_sfixed(-0.9422,1,L_SIZE),
				to_sfixed(-0.9421,1,L_SIZE),
				to_sfixed(-0.9421,1,L_SIZE),
				to_sfixed(-0.9421,1,L_SIZE),
				to_sfixed(-0.9420,1,L_SIZE),
				to_sfixed(-0.9420,1,L_SIZE),
				to_sfixed(-0.9419,1,L_SIZE),
				to_sfixed(-0.9419,1,L_SIZE),
				to_sfixed(-0.9418,1,L_SIZE),
				to_sfixed(-0.9418,1,L_SIZE),
				to_sfixed(-0.9418,1,L_SIZE),
				to_sfixed(-0.9417,1,L_SIZE),
				to_sfixed(-0.9417,1,L_SIZE),
				to_sfixed(-0.9416,1,L_SIZE),
				to_sfixed(-0.9416,1,L_SIZE),
				to_sfixed(-0.9416,1,L_SIZE),
				to_sfixed(-0.9415,1,L_SIZE),
				to_sfixed(-0.9415,1,L_SIZE),
				to_sfixed(-0.9414,1,L_SIZE),
				to_sfixed(-0.9414,1,L_SIZE),
				to_sfixed(-0.9413,1,L_SIZE),
				to_sfixed(-0.9413,1,L_SIZE),
				to_sfixed(-0.9413,1,L_SIZE),
				to_sfixed(-0.9412,1,L_SIZE),
				to_sfixed(-0.9412,1,L_SIZE),
				to_sfixed(-0.9411,1,L_SIZE),
				to_sfixed(-0.9411,1,L_SIZE),
				to_sfixed(-0.9411,1,L_SIZE),
				to_sfixed(-0.9410,1,L_SIZE),
				to_sfixed(-0.9410,1,L_SIZE),
				to_sfixed(-0.9409,1,L_SIZE),
				to_sfixed(-0.9409,1,L_SIZE),
				to_sfixed(-0.9408,1,L_SIZE),
				to_sfixed(-0.9408,1,L_SIZE),
				to_sfixed(-0.9408,1,L_SIZE),
				to_sfixed(-0.9407,1,L_SIZE),
				to_sfixed(-0.9407,1,L_SIZE),
				to_sfixed(-0.9406,1,L_SIZE),
				to_sfixed(-0.9406,1,L_SIZE),
				to_sfixed(-0.9406,1,L_SIZE),
				to_sfixed(-0.9405,1,L_SIZE),
				to_sfixed(-0.9405,1,L_SIZE),
				to_sfixed(-0.9404,1,L_SIZE),
				to_sfixed(-0.9404,1,L_SIZE),
				to_sfixed(-0.9403,1,L_SIZE),
				to_sfixed(-0.9403,1,L_SIZE),
				to_sfixed(-0.9403,1,L_SIZE),
				to_sfixed(-0.9402,1,L_SIZE),
				to_sfixed(-0.9402,1,L_SIZE),
				to_sfixed(-0.9401,1,L_SIZE),
				to_sfixed(-0.9401,1,L_SIZE),
				to_sfixed(-0.9400,1,L_SIZE),
				to_sfixed(-0.9400,1,L_SIZE),
				to_sfixed(-0.9400,1,L_SIZE),
				to_sfixed(-0.9399,1,L_SIZE),
				to_sfixed(-0.9399,1,L_SIZE),
				to_sfixed(-0.9398,1,L_SIZE),
				to_sfixed(-0.9398,1,L_SIZE),
				to_sfixed(-0.9397,1,L_SIZE),
				to_sfixed(-0.9397,1,L_SIZE),
				to_sfixed(-0.9397,1,L_SIZE),
				to_sfixed(-0.9396,1,L_SIZE),
				to_sfixed(-0.9396,1,L_SIZE),
				to_sfixed(-0.9395,1,L_SIZE),
				to_sfixed(-0.9395,1,L_SIZE),
				to_sfixed(-0.9394,1,L_SIZE),
				to_sfixed(-0.9394,1,L_SIZE),
				to_sfixed(-0.9394,1,L_SIZE),
				to_sfixed(-0.9393,1,L_SIZE),
				to_sfixed(-0.9393,1,L_SIZE),
				to_sfixed(-0.9392,1,L_SIZE),
				to_sfixed(-0.9392,1,L_SIZE),
				to_sfixed(-0.9391,1,L_SIZE),
				to_sfixed(-0.9391,1,L_SIZE),
				to_sfixed(-0.9391,1,L_SIZE),
				to_sfixed(-0.9390,1,L_SIZE),
				to_sfixed(-0.9390,1,L_SIZE),
				to_sfixed(-0.9389,1,L_SIZE),
				to_sfixed(-0.9389,1,L_SIZE),
				to_sfixed(-0.9388,1,L_SIZE),
				to_sfixed(-0.9388,1,L_SIZE),
				to_sfixed(-0.9387,1,L_SIZE),
				to_sfixed(-0.9387,1,L_SIZE),
				to_sfixed(-0.9387,1,L_SIZE),
				to_sfixed(-0.9386,1,L_SIZE),
				to_sfixed(-0.9386,1,L_SIZE),
				to_sfixed(-0.9385,1,L_SIZE),
				to_sfixed(-0.9385,1,L_SIZE),
				to_sfixed(-0.9384,1,L_SIZE),
				to_sfixed(-0.9384,1,L_SIZE),
				to_sfixed(-0.9384,1,L_SIZE),
				to_sfixed(-0.9383,1,L_SIZE),
				to_sfixed(-0.9383,1,L_SIZE),
				to_sfixed(-0.9382,1,L_SIZE),
				to_sfixed(-0.9382,1,L_SIZE),
				to_sfixed(-0.9381,1,L_SIZE),
				to_sfixed(-0.9381,1,L_SIZE),
				to_sfixed(-0.9381,1,L_SIZE),
				to_sfixed(-0.9380,1,L_SIZE),
				to_sfixed(-0.9380,1,L_SIZE),
				to_sfixed(-0.9379,1,L_SIZE),
				to_sfixed(-0.9379,1,L_SIZE),
				to_sfixed(-0.9378,1,L_SIZE),
				to_sfixed(-0.9378,1,L_SIZE),
				to_sfixed(-0.9377,1,L_SIZE),
				to_sfixed(-0.9377,1,L_SIZE),
				to_sfixed(-0.9377,1,L_SIZE),
				to_sfixed(-0.9376,1,L_SIZE),
				to_sfixed(-0.9376,1,L_SIZE),
				to_sfixed(-0.9375,1,L_SIZE),
				to_sfixed(-0.9375,1,L_SIZE),
				to_sfixed(-0.9374,1,L_SIZE),
				to_sfixed(-0.9374,1,L_SIZE),
				to_sfixed(-0.9373,1,L_SIZE),
				to_sfixed(-0.9373,1,L_SIZE),
				to_sfixed(-0.9373,1,L_SIZE),
				to_sfixed(-0.9372,1,L_SIZE),
				to_sfixed(-0.9372,1,L_SIZE),
				to_sfixed(-0.9371,1,L_SIZE),
				to_sfixed(-0.9371,1,L_SIZE),
				to_sfixed(-0.9370,1,L_SIZE),
				to_sfixed(-0.9370,1,L_SIZE),
				to_sfixed(-0.9369,1,L_SIZE),
				to_sfixed(-0.9369,1,L_SIZE),
				to_sfixed(-0.9369,1,L_SIZE),
				to_sfixed(-0.9368,1,L_SIZE),
				to_sfixed(-0.9368,1,L_SIZE),
				to_sfixed(-0.9367,1,L_SIZE),
				to_sfixed(-0.9367,1,L_SIZE),
				to_sfixed(-0.9366,1,L_SIZE),
				to_sfixed(-0.9366,1,L_SIZE),
				to_sfixed(-0.9365,1,L_SIZE),
				to_sfixed(-0.9365,1,L_SIZE),
				to_sfixed(-0.9364,1,L_SIZE),
				to_sfixed(-0.9364,1,L_SIZE),
				to_sfixed(-0.9364,1,L_SIZE),
				to_sfixed(-0.9363,1,L_SIZE),
				to_sfixed(-0.9363,1,L_SIZE),
				to_sfixed(-0.9362,1,L_SIZE),
				to_sfixed(-0.9362,1,L_SIZE),
				to_sfixed(-0.9361,1,L_SIZE),
				to_sfixed(-0.9361,1,L_SIZE),
				to_sfixed(-0.9360,1,L_SIZE),
				to_sfixed(-0.9360,1,L_SIZE),
				to_sfixed(-0.9360,1,L_SIZE),
				to_sfixed(-0.9359,1,L_SIZE),
				to_sfixed(-0.9359,1,L_SIZE),
				to_sfixed(-0.9358,1,L_SIZE),
				to_sfixed(-0.9358,1,L_SIZE),
				to_sfixed(-0.9357,1,L_SIZE),
				to_sfixed(-0.9357,1,L_SIZE),
				to_sfixed(-0.9356,1,L_SIZE),
				to_sfixed(-0.9356,1,L_SIZE),
				to_sfixed(-0.9355,1,L_SIZE),
				to_sfixed(-0.9355,1,L_SIZE),
				to_sfixed(-0.9354,1,L_SIZE),
				to_sfixed(-0.9354,1,L_SIZE),
				to_sfixed(-0.9354,1,L_SIZE),
				to_sfixed(-0.9353,1,L_SIZE),
				to_sfixed(-0.9353,1,L_SIZE),
				to_sfixed(-0.9352,1,L_SIZE),
				to_sfixed(-0.9352,1,L_SIZE),
				to_sfixed(-0.9351,1,L_SIZE),
				to_sfixed(-0.9351,1,L_SIZE),
				to_sfixed(-0.9350,1,L_SIZE),
				to_sfixed(-0.9350,1,L_SIZE),
				to_sfixed(-0.9349,1,L_SIZE),
				to_sfixed(-0.9349,1,L_SIZE),
				to_sfixed(-0.9349,1,L_SIZE),
				to_sfixed(-0.9348,1,L_SIZE),
				to_sfixed(-0.9348,1,L_SIZE),
				to_sfixed(-0.9347,1,L_SIZE),
				to_sfixed(-0.9347,1,L_SIZE),
				to_sfixed(-0.9346,1,L_SIZE),
				to_sfixed(-0.9346,1,L_SIZE),
				to_sfixed(-0.9345,1,L_SIZE),
				to_sfixed(-0.9345,1,L_SIZE),
				to_sfixed(-0.9344,1,L_SIZE),
				to_sfixed(-0.9344,1,L_SIZE),
				to_sfixed(-0.9343,1,L_SIZE),
				to_sfixed(-0.9343,1,L_SIZE),
				to_sfixed(-0.9342,1,L_SIZE),
				to_sfixed(-0.9342,1,L_SIZE),
				to_sfixed(-0.9342,1,L_SIZE),
				to_sfixed(-0.9341,1,L_SIZE),
				to_sfixed(-0.9341,1,L_SIZE),
				to_sfixed(-0.9340,1,L_SIZE),
				to_sfixed(-0.9340,1,L_SIZE),
				to_sfixed(-0.9339,1,L_SIZE),
				to_sfixed(-0.9339,1,L_SIZE),
				to_sfixed(-0.9338,1,L_SIZE),
				to_sfixed(-0.9338,1,L_SIZE),
				to_sfixed(-0.9337,1,L_SIZE),
				to_sfixed(-0.9337,1,L_SIZE),
				to_sfixed(-0.9336,1,L_SIZE),
				to_sfixed(-0.9336,1,L_SIZE),
				to_sfixed(-0.9335,1,L_SIZE),
				to_sfixed(-0.9335,1,L_SIZE),
				to_sfixed(-0.9335,1,L_SIZE),
				to_sfixed(-0.9334,1,L_SIZE),
				to_sfixed(-0.9334,1,L_SIZE),
				to_sfixed(-0.9333,1,L_SIZE),
				to_sfixed(-0.9333,1,L_SIZE),
				to_sfixed(-0.9332,1,L_SIZE),
				to_sfixed(-0.9332,1,L_SIZE),
				to_sfixed(-0.9331,1,L_SIZE),
				to_sfixed(-0.9331,1,L_SIZE),
				to_sfixed(-0.9330,1,L_SIZE),
				to_sfixed(-0.9330,1,L_SIZE),
				to_sfixed(-0.9329,1,L_SIZE),
				to_sfixed(-0.9329,1,L_SIZE),
				to_sfixed(-0.9328,1,L_SIZE),
				to_sfixed(-0.9328,1,L_SIZE),
				to_sfixed(-0.9327,1,L_SIZE),
				to_sfixed(-0.9327,1,L_SIZE),
				to_sfixed(-0.9326,1,L_SIZE),
				to_sfixed(-0.9326,1,L_SIZE),
				to_sfixed(-0.9326,1,L_SIZE),
				to_sfixed(-0.9325,1,L_SIZE),
				to_sfixed(-0.9325,1,L_SIZE),
				to_sfixed(-0.9324,1,L_SIZE),
				to_sfixed(-0.9324,1,L_SIZE),
				to_sfixed(-0.9323,1,L_SIZE),
				to_sfixed(-0.9323,1,L_SIZE),
				to_sfixed(-0.9322,1,L_SIZE),
				to_sfixed(-0.9322,1,L_SIZE),
				to_sfixed(-0.9321,1,L_SIZE),
				to_sfixed(-0.9321,1,L_SIZE),
				to_sfixed(-0.9320,1,L_SIZE),
				to_sfixed(-0.9320,1,L_SIZE),
				to_sfixed(-0.9319,1,L_SIZE),
				to_sfixed(-0.9319,1,L_SIZE),
				to_sfixed(-0.9318,1,L_SIZE),
				to_sfixed(-0.9318,1,L_SIZE),
				to_sfixed(-0.9317,1,L_SIZE),
				to_sfixed(-0.9317,1,L_SIZE),
				to_sfixed(-0.9316,1,L_SIZE),
				to_sfixed(-0.9316,1,L_SIZE),
				to_sfixed(-0.9315,1,L_SIZE),
				to_sfixed(-0.9315,1,L_SIZE),
				to_sfixed(-0.9314,1,L_SIZE),
				to_sfixed(-0.9314,1,L_SIZE),
				to_sfixed(-0.9313,1,L_SIZE),
				to_sfixed(-0.9313,1,L_SIZE),
				to_sfixed(-0.9313,1,L_SIZE),
				to_sfixed(-0.9312,1,L_SIZE),
				to_sfixed(-0.9312,1,L_SIZE),
				to_sfixed(-0.9311,1,L_SIZE),
				to_sfixed(-0.9311,1,L_SIZE),
				to_sfixed(-0.9310,1,L_SIZE),
				to_sfixed(-0.9310,1,L_SIZE),
				to_sfixed(-0.9309,1,L_SIZE),
				to_sfixed(-0.9309,1,L_SIZE),
				to_sfixed(-0.9308,1,L_SIZE),
				to_sfixed(-0.9308,1,L_SIZE),
				to_sfixed(-0.9307,1,L_SIZE),
				to_sfixed(-0.9307,1,L_SIZE),
				to_sfixed(-0.9306,1,L_SIZE),
				to_sfixed(-0.9306,1,L_SIZE),
				to_sfixed(-0.9305,1,L_SIZE),
				to_sfixed(-0.9305,1,L_SIZE),
				to_sfixed(-0.9304,1,L_SIZE),
				to_sfixed(-0.9304,1,L_SIZE),
				to_sfixed(-0.9303,1,L_SIZE),
				to_sfixed(-0.9303,1,L_SIZE),
				to_sfixed(-0.9302,1,L_SIZE),
				to_sfixed(-0.9302,1,L_SIZE),
				to_sfixed(-0.9301,1,L_SIZE),
				to_sfixed(-0.9301,1,L_SIZE),
				to_sfixed(-0.9300,1,L_SIZE),
				to_sfixed(-0.9300,1,L_SIZE),
				to_sfixed(-0.9299,1,L_SIZE),
				to_sfixed(-0.9299,1,L_SIZE),
				to_sfixed(-0.9298,1,L_SIZE),
				to_sfixed(-0.9298,1,L_SIZE),
				to_sfixed(-0.9297,1,L_SIZE),
				to_sfixed(-0.9297,1,L_SIZE),
				to_sfixed(-0.9296,1,L_SIZE),
				to_sfixed(-0.9296,1,L_SIZE),
				to_sfixed(-0.9295,1,L_SIZE),
				to_sfixed(-0.9295,1,L_SIZE),
				to_sfixed(-0.9294,1,L_SIZE),
				to_sfixed(-0.9294,1,L_SIZE),
				to_sfixed(-0.9293,1,L_SIZE),
				to_sfixed(-0.9293,1,L_SIZE),
				to_sfixed(-0.9292,1,L_SIZE),
				to_sfixed(-0.9292,1,L_SIZE),
				to_sfixed(-0.9291,1,L_SIZE),
				to_sfixed(-0.9291,1,L_SIZE),
				to_sfixed(-0.9290,1,L_SIZE),
				to_sfixed(-0.9290,1,L_SIZE),
				to_sfixed(-0.9289,1,L_SIZE),
				to_sfixed(-0.9289,1,L_SIZE),
				to_sfixed(-0.9288,1,L_SIZE),
				to_sfixed(-0.9288,1,L_SIZE),
				to_sfixed(-0.9287,1,L_SIZE),
				to_sfixed(-0.9287,1,L_SIZE),
				to_sfixed(-0.9286,1,L_SIZE),
				to_sfixed(-0.9286,1,L_SIZE),
				to_sfixed(-0.9285,1,L_SIZE),
				to_sfixed(-0.9285,1,L_SIZE),
				to_sfixed(-0.9284,1,L_SIZE),
				to_sfixed(-0.9284,1,L_SIZE),
				to_sfixed(-0.9283,1,L_SIZE),
				to_sfixed(-0.9283,1,L_SIZE),
				to_sfixed(-0.9282,1,L_SIZE),
				to_sfixed(-0.9282,1,L_SIZE),
				to_sfixed(-0.9281,1,L_SIZE),
				to_sfixed(-0.9281,1,L_SIZE),
				to_sfixed(-0.9280,1,L_SIZE),
				to_sfixed(-0.9280,1,L_SIZE),
				to_sfixed(-0.9279,1,L_SIZE),
				to_sfixed(-0.9279,1,L_SIZE),
				to_sfixed(-0.9278,1,L_SIZE),
				to_sfixed(-0.9278,1,L_SIZE),
				to_sfixed(-0.9277,1,L_SIZE),
				to_sfixed(-0.9277,1,L_SIZE),
				to_sfixed(-0.9276,1,L_SIZE),
				to_sfixed(-0.9276,1,L_SIZE),
				to_sfixed(-0.9275,1,L_SIZE),
				to_sfixed(-0.9275,1,L_SIZE),
				to_sfixed(-0.9274,1,L_SIZE),
				to_sfixed(-0.9274,1,L_SIZE),
				to_sfixed(-0.9273,1,L_SIZE),
				to_sfixed(-0.9273,1,L_SIZE),
				to_sfixed(-0.9272,1,L_SIZE),
				to_sfixed(-0.9271,1,L_SIZE),
				to_sfixed(-0.9271,1,L_SIZE),
				to_sfixed(-0.9270,1,L_SIZE),
				to_sfixed(-0.9270,1,L_SIZE),
				to_sfixed(-0.9269,1,L_SIZE),
				to_sfixed(-0.9269,1,L_SIZE),
				to_sfixed(-0.9268,1,L_SIZE),
				to_sfixed(-0.9268,1,L_SIZE),
				to_sfixed(-0.9267,1,L_SIZE),
				to_sfixed(-0.9267,1,L_SIZE),
				to_sfixed(-0.9266,1,L_SIZE),
				to_sfixed(-0.9266,1,L_SIZE),
				to_sfixed(-0.9265,1,L_SIZE),
				to_sfixed(-0.9265,1,L_SIZE),
				to_sfixed(-0.9264,1,L_SIZE),
				to_sfixed(-0.9264,1,L_SIZE),
				to_sfixed(-0.9263,1,L_SIZE),
				to_sfixed(-0.9263,1,L_SIZE),
				to_sfixed(-0.9262,1,L_SIZE),
				to_sfixed(-0.9262,1,L_SIZE),
				to_sfixed(-0.9261,1,L_SIZE),
				to_sfixed(-0.9261,1,L_SIZE),
				to_sfixed(-0.9260,1,L_SIZE),
				to_sfixed(-0.9260,1,L_SIZE),
				to_sfixed(-0.9259,1,L_SIZE),
				to_sfixed(-0.9259,1,L_SIZE),
				to_sfixed(-0.9258,1,L_SIZE),
				to_sfixed(-0.9257,1,L_SIZE),
				to_sfixed(-0.9257,1,L_SIZE),
				to_sfixed(-0.9256,1,L_SIZE),
				to_sfixed(-0.9256,1,L_SIZE),
				to_sfixed(-0.9255,1,L_SIZE),
				to_sfixed(-0.9255,1,L_SIZE),
				to_sfixed(-0.9254,1,L_SIZE),
				to_sfixed(-0.9254,1,L_SIZE),
				to_sfixed(-0.9253,1,L_SIZE),
				to_sfixed(-0.9253,1,L_SIZE),
				to_sfixed(-0.9252,1,L_SIZE),
				to_sfixed(-0.9252,1,L_SIZE),
				to_sfixed(-0.9251,1,L_SIZE),
				to_sfixed(-0.9251,1,L_SIZE),
				to_sfixed(-0.9250,1,L_SIZE),
				to_sfixed(-0.9250,1,L_SIZE),
				to_sfixed(-0.9249,1,L_SIZE),
				to_sfixed(-0.9249,1,L_SIZE),
				to_sfixed(-0.9248,1,L_SIZE),
				to_sfixed(-0.9247,1,L_SIZE),
				to_sfixed(-0.9247,1,L_SIZE),
				to_sfixed(-0.9246,1,L_SIZE),
				to_sfixed(-0.9246,1,L_SIZE),
				to_sfixed(-0.9245,1,L_SIZE),
				to_sfixed(-0.9245,1,L_SIZE),
				to_sfixed(-0.9244,1,L_SIZE),
				to_sfixed(-0.9244,1,L_SIZE),
				to_sfixed(-0.9243,1,L_SIZE),
				to_sfixed(-0.9243,1,L_SIZE),
				to_sfixed(-0.9242,1,L_SIZE),
				to_sfixed(-0.9242,1,L_SIZE),
				to_sfixed(-0.9241,1,L_SIZE),
				to_sfixed(-0.9241,1,L_SIZE),
				to_sfixed(-0.9240,1,L_SIZE),
				to_sfixed(-0.9239,1,L_SIZE),
				to_sfixed(-0.9239,1,L_SIZE),
				to_sfixed(-0.9238,1,L_SIZE),
				to_sfixed(-0.9238,1,L_SIZE),
				to_sfixed(-0.9237,1,L_SIZE),
				to_sfixed(-0.9237,1,L_SIZE),
				to_sfixed(-0.9236,1,L_SIZE),
				to_sfixed(-0.9236,1,L_SIZE),
				to_sfixed(-0.9235,1,L_SIZE),
				to_sfixed(-0.9235,1,L_SIZE),
				to_sfixed(-0.9234,1,L_SIZE),
				to_sfixed(-0.9234,1,L_SIZE),
				to_sfixed(-0.9233,1,L_SIZE),
				to_sfixed(-0.9232,1,L_SIZE),
				to_sfixed(-0.9232,1,L_SIZE),
				to_sfixed(-0.9231,1,L_SIZE),
				to_sfixed(-0.9231,1,L_SIZE),
				to_sfixed(-0.9230,1,L_SIZE),
				to_sfixed(-0.9230,1,L_SIZE),
				to_sfixed(-0.9229,1,L_SIZE),
				to_sfixed(-0.9229,1,L_SIZE),
				to_sfixed(-0.9228,1,L_SIZE),
				to_sfixed(-0.9228,1,L_SIZE),
				to_sfixed(-0.9227,1,L_SIZE),
				to_sfixed(-0.9227,1,L_SIZE),
				to_sfixed(-0.9226,1,L_SIZE),
				to_sfixed(-0.9225,1,L_SIZE),
				to_sfixed(-0.9225,1,L_SIZE),
				to_sfixed(-0.9224,1,L_SIZE),
				to_sfixed(-0.9224,1,L_SIZE),
				to_sfixed(-0.9223,1,L_SIZE),
				to_sfixed(-0.9223,1,L_SIZE),
				to_sfixed(-0.9222,1,L_SIZE),
				to_sfixed(-0.9222,1,L_SIZE),
				to_sfixed(-0.9221,1,L_SIZE),
				to_sfixed(-0.9220,1,L_SIZE),
				to_sfixed(-0.9220,1,L_SIZE),
				to_sfixed(-0.9219,1,L_SIZE),
				to_sfixed(-0.9219,1,L_SIZE),
				to_sfixed(-0.9218,1,L_SIZE),
				to_sfixed(-0.9218,1,L_SIZE),
				to_sfixed(-0.9217,1,L_SIZE),
				to_sfixed(-0.9217,1,L_SIZE),
				to_sfixed(-0.9216,1,L_SIZE),
				to_sfixed(-0.9216,1,L_SIZE),
				to_sfixed(-0.9215,1,L_SIZE),
				to_sfixed(-0.9214,1,L_SIZE),
				to_sfixed(-0.9214,1,L_SIZE),
				to_sfixed(-0.9213,1,L_SIZE),
				to_sfixed(-0.9213,1,L_SIZE),
				to_sfixed(-0.9212,1,L_SIZE),
				to_sfixed(-0.9212,1,L_SIZE),
				to_sfixed(-0.9211,1,L_SIZE),
				to_sfixed(-0.9211,1,L_SIZE),
				to_sfixed(-0.9210,1,L_SIZE),
				to_sfixed(-0.9209,1,L_SIZE),
				to_sfixed(-0.9209,1,L_SIZE),
				to_sfixed(-0.9208,1,L_SIZE),
				to_sfixed(-0.9208,1,L_SIZE),
				to_sfixed(-0.9207,1,L_SIZE),
				to_sfixed(-0.9207,1,L_SIZE),
				to_sfixed(-0.9206,1,L_SIZE),
				to_sfixed(-0.9206,1,L_SIZE),
				to_sfixed(-0.9205,1,L_SIZE),
				to_sfixed(-0.9204,1,L_SIZE),
				to_sfixed(-0.9204,1,L_SIZE),
				to_sfixed(-0.9203,1,L_SIZE),
				to_sfixed(-0.9203,1,L_SIZE),
				to_sfixed(-0.9202,1,L_SIZE),
				to_sfixed(-0.9202,1,L_SIZE),
				to_sfixed(-0.9201,1,L_SIZE),
				to_sfixed(-0.9201,1,L_SIZE),
				to_sfixed(-0.9200,1,L_SIZE),
				to_sfixed(-0.9199,1,L_SIZE),
				to_sfixed(-0.9199,1,L_SIZE),
				to_sfixed(-0.9198,1,L_SIZE),
				to_sfixed(-0.9198,1,L_SIZE),
				to_sfixed(-0.9197,1,L_SIZE),
				to_sfixed(-0.9197,1,L_SIZE),
				to_sfixed(-0.9196,1,L_SIZE),
				to_sfixed(-0.9195,1,L_SIZE),
				to_sfixed(-0.9195,1,L_SIZE),
				to_sfixed(-0.9194,1,L_SIZE),
				to_sfixed(-0.9194,1,L_SIZE),
				to_sfixed(-0.9193,1,L_SIZE),
				to_sfixed(-0.9193,1,L_SIZE),
				to_sfixed(-0.9192,1,L_SIZE),
				to_sfixed(-0.9191,1,L_SIZE),
				to_sfixed(-0.9191,1,L_SIZE),
				to_sfixed(-0.9190,1,L_SIZE),
				to_sfixed(-0.9190,1,L_SIZE),
				to_sfixed(-0.9189,1,L_SIZE),
				to_sfixed(-0.9189,1,L_SIZE),
				to_sfixed(-0.9188,1,L_SIZE),
				to_sfixed(-0.9187,1,L_SIZE),
				to_sfixed(-0.9187,1,L_SIZE),
				to_sfixed(-0.9186,1,L_SIZE),
				to_sfixed(-0.9186,1,L_SIZE),
				to_sfixed(-0.9185,1,L_SIZE),
				to_sfixed(-0.9185,1,L_SIZE),
				to_sfixed(-0.9184,1,L_SIZE),
				to_sfixed(-0.9183,1,L_SIZE),
				to_sfixed(-0.9183,1,L_SIZE),
				to_sfixed(-0.9182,1,L_SIZE),
				to_sfixed(-0.9182,1,L_SIZE),
				to_sfixed(-0.9181,1,L_SIZE),
				to_sfixed(-0.9181,1,L_SIZE),
				to_sfixed(-0.9180,1,L_SIZE),
				to_sfixed(-0.9179,1,L_SIZE),
				to_sfixed(-0.9179,1,L_SIZE),
				to_sfixed(-0.9178,1,L_SIZE),
				to_sfixed(-0.9178,1,L_SIZE),
				to_sfixed(-0.9177,1,L_SIZE),
				to_sfixed(-0.9177,1,L_SIZE),
				to_sfixed(-0.9176,1,L_SIZE),
				to_sfixed(-0.9175,1,L_SIZE),
				to_sfixed(-0.9175,1,L_SIZE),
				to_sfixed(-0.9174,1,L_SIZE),
				to_sfixed(-0.9174,1,L_SIZE),
				to_sfixed(-0.9173,1,L_SIZE),
				to_sfixed(-0.9172,1,L_SIZE),
				to_sfixed(-0.9172,1,L_SIZE),
				to_sfixed(-0.9171,1,L_SIZE),
				to_sfixed(-0.9171,1,L_SIZE),
				to_sfixed(-0.9170,1,L_SIZE),
				to_sfixed(-0.9170,1,L_SIZE),
				to_sfixed(-0.9169,1,L_SIZE),
				to_sfixed(-0.9168,1,L_SIZE),
				to_sfixed(-0.9168,1,L_SIZE),
				to_sfixed(-0.9167,1,L_SIZE),
				to_sfixed(-0.9167,1,L_SIZE),
				to_sfixed(-0.9166,1,L_SIZE),
				to_sfixed(-0.9165,1,L_SIZE),
				to_sfixed(-0.9165,1,L_SIZE),
				to_sfixed(-0.9164,1,L_SIZE),
				to_sfixed(-0.9164,1,L_SIZE),
				to_sfixed(-0.9163,1,L_SIZE),
				to_sfixed(-0.9163,1,L_SIZE),
				to_sfixed(-0.9162,1,L_SIZE),
				to_sfixed(-0.9161,1,L_SIZE),
				to_sfixed(-0.9161,1,L_SIZE),
				to_sfixed(-0.9160,1,L_SIZE),
				to_sfixed(-0.9160,1,L_SIZE),
				to_sfixed(-0.9159,1,L_SIZE),
				to_sfixed(-0.9158,1,L_SIZE),
				to_sfixed(-0.9158,1,L_SIZE),
				to_sfixed(-0.9157,1,L_SIZE),
				to_sfixed(-0.9157,1,L_SIZE),
				to_sfixed(-0.9156,1,L_SIZE),
				to_sfixed(-0.9155,1,L_SIZE),
				to_sfixed(-0.9155,1,L_SIZE),
				to_sfixed(-0.9154,1,L_SIZE),
				to_sfixed(-0.9154,1,L_SIZE),
				to_sfixed(-0.9153,1,L_SIZE),
				to_sfixed(-0.9153,1,L_SIZE),
				to_sfixed(-0.9152,1,L_SIZE),
				to_sfixed(-0.9151,1,L_SIZE),
				to_sfixed(-0.9151,1,L_SIZE),
				to_sfixed(-0.9150,1,L_SIZE),
				to_sfixed(-0.9150,1,L_SIZE),
				to_sfixed(-0.9149,1,L_SIZE),
				to_sfixed(-0.9148,1,L_SIZE),
				to_sfixed(-0.9148,1,L_SIZE),
				to_sfixed(-0.9147,1,L_SIZE),
				to_sfixed(-0.9147,1,L_SIZE),
				to_sfixed(-0.9146,1,L_SIZE),
				to_sfixed(-0.9145,1,L_SIZE),
				to_sfixed(-0.9145,1,L_SIZE),
				to_sfixed(-0.9144,1,L_SIZE),
				to_sfixed(-0.9144,1,L_SIZE),
				to_sfixed(-0.9143,1,L_SIZE),
				to_sfixed(-0.9142,1,L_SIZE),
				to_sfixed(-0.9142,1,L_SIZE),
				to_sfixed(-0.9141,1,L_SIZE),
				to_sfixed(-0.9141,1,L_SIZE),
				to_sfixed(-0.9140,1,L_SIZE),
				to_sfixed(-0.9139,1,L_SIZE),
				to_sfixed(-0.9139,1,L_SIZE),
				to_sfixed(-0.9138,1,L_SIZE),
				to_sfixed(-0.9138,1,L_SIZE),
				to_sfixed(-0.9137,1,L_SIZE),
				to_sfixed(-0.9136,1,L_SIZE),
				to_sfixed(-0.9136,1,L_SIZE),
				to_sfixed(-0.9135,1,L_SIZE),
				to_sfixed(-0.9135,1,L_SIZE),
				to_sfixed(-0.9134,1,L_SIZE),
				to_sfixed(-0.9133,1,L_SIZE),
				to_sfixed(-0.9133,1,L_SIZE),
				to_sfixed(-0.9132,1,L_SIZE),
				to_sfixed(-0.9131,1,L_SIZE),
				to_sfixed(-0.9131,1,L_SIZE),
				to_sfixed(-0.9130,1,L_SIZE),
				to_sfixed(-0.9130,1,L_SIZE),
				to_sfixed(-0.9129,1,L_SIZE),
				to_sfixed(-0.9128,1,L_SIZE),
				to_sfixed(-0.9128,1,L_SIZE),
				to_sfixed(-0.9127,1,L_SIZE),
				to_sfixed(-0.9127,1,L_SIZE),
				to_sfixed(-0.9126,1,L_SIZE),
				to_sfixed(-0.9125,1,L_SIZE),
				to_sfixed(-0.9125,1,L_SIZE),
				to_sfixed(-0.9124,1,L_SIZE),
				to_sfixed(-0.9124,1,L_SIZE),
				to_sfixed(-0.9123,1,L_SIZE),
				to_sfixed(-0.9122,1,L_SIZE),
				to_sfixed(-0.9122,1,L_SIZE),
				to_sfixed(-0.9121,1,L_SIZE),
				to_sfixed(-0.9120,1,L_SIZE),
				to_sfixed(-0.9120,1,L_SIZE),
				to_sfixed(-0.9119,1,L_SIZE),
				to_sfixed(-0.9119,1,L_SIZE),
				to_sfixed(-0.9118,1,L_SIZE),
				to_sfixed(-0.9117,1,L_SIZE),
				to_sfixed(-0.9117,1,L_SIZE),
				to_sfixed(-0.9116,1,L_SIZE),
				to_sfixed(-0.9116,1,L_SIZE),
				to_sfixed(-0.9115,1,L_SIZE),
				to_sfixed(-0.9114,1,L_SIZE),
				to_sfixed(-0.9114,1,L_SIZE),
				to_sfixed(-0.9113,1,L_SIZE),
				to_sfixed(-0.9112,1,L_SIZE),
				to_sfixed(-0.9112,1,L_SIZE),
				to_sfixed(-0.9111,1,L_SIZE),
				to_sfixed(-0.9111,1,L_SIZE),
				to_sfixed(-0.9110,1,L_SIZE),
				to_sfixed(-0.9109,1,L_SIZE),
				to_sfixed(-0.9109,1,L_SIZE),
				to_sfixed(-0.9108,1,L_SIZE),
				to_sfixed(-0.9107,1,L_SIZE),
				to_sfixed(-0.9107,1,L_SIZE),
				to_sfixed(-0.9106,1,L_SIZE),
				to_sfixed(-0.9106,1,L_SIZE),
				to_sfixed(-0.9105,1,L_SIZE),
				to_sfixed(-0.9104,1,L_SIZE),
				to_sfixed(-0.9104,1,L_SIZE),
				to_sfixed(-0.9103,1,L_SIZE),
				to_sfixed(-0.9102,1,L_SIZE),
				to_sfixed(-0.9102,1,L_SIZE),
				to_sfixed(-0.9101,1,L_SIZE),
				to_sfixed(-0.9101,1,L_SIZE),
				to_sfixed(-0.9100,1,L_SIZE),
				to_sfixed(-0.9099,1,L_SIZE),
				to_sfixed(-0.9099,1,L_SIZE),
				to_sfixed(-0.9098,1,L_SIZE),
				to_sfixed(-0.9097,1,L_SIZE),
				to_sfixed(-0.9097,1,L_SIZE),
				to_sfixed(-0.9096,1,L_SIZE),
				to_sfixed(-0.9095,1,L_SIZE),
				to_sfixed(-0.9095,1,L_SIZE),
				to_sfixed(-0.9094,1,L_SIZE),
				to_sfixed(-0.9094,1,L_SIZE),
				to_sfixed(-0.9093,1,L_SIZE),
				to_sfixed(-0.9092,1,L_SIZE),
				to_sfixed(-0.9092,1,L_SIZE),
				to_sfixed(-0.9091,1,L_SIZE),
				to_sfixed(-0.9090,1,L_SIZE),
				to_sfixed(-0.9090,1,L_SIZE),
				to_sfixed(-0.9089,1,L_SIZE),
				to_sfixed(-0.9088,1,L_SIZE),
				to_sfixed(-0.9088,1,L_SIZE),
				to_sfixed(-0.9087,1,L_SIZE),
				to_sfixed(-0.9087,1,L_SIZE),
				to_sfixed(-0.9086,1,L_SIZE),
				to_sfixed(-0.9085,1,L_SIZE),
				to_sfixed(-0.9085,1,L_SIZE),
				to_sfixed(-0.9084,1,L_SIZE),
				to_sfixed(-0.9083,1,L_SIZE),
				to_sfixed(-0.9083,1,L_SIZE),
				to_sfixed(-0.9082,1,L_SIZE),
				to_sfixed(-0.9081,1,L_SIZE),
				to_sfixed(-0.9081,1,L_SIZE),
				to_sfixed(-0.9080,1,L_SIZE),
				to_sfixed(-0.9080,1,L_SIZE),
				to_sfixed(-0.9079,1,L_SIZE),
				to_sfixed(-0.9078,1,L_SIZE),
				to_sfixed(-0.9078,1,L_SIZE),
				to_sfixed(-0.9077,1,L_SIZE),
				to_sfixed(-0.9076,1,L_SIZE),
				to_sfixed(-0.9076,1,L_SIZE),
				to_sfixed(-0.9075,1,L_SIZE),
				to_sfixed(-0.9074,1,L_SIZE),
				to_sfixed(-0.9074,1,L_SIZE),
				to_sfixed(-0.9073,1,L_SIZE),
				to_sfixed(-0.9072,1,L_SIZE),
				to_sfixed(-0.9072,1,L_SIZE),
				to_sfixed(-0.9071,1,L_SIZE),
				to_sfixed(-0.9070,1,L_SIZE),
				to_sfixed(-0.9070,1,L_SIZE),
				to_sfixed(-0.9069,1,L_SIZE),
				to_sfixed(-0.9069,1,L_SIZE),
				to_sfixed(-0.9068,1,L_SIZE),
				to_sfixed(-0.9067,1,L_SIZE),
				to_sfixed(-0.9067,1,L_SIZE),
				to_sfixed(-0.9066,1,L_SIZE),
				to_sfixed(-0.9065,1,L_SIZE),
				to_sfixed(-0.9065,1,L_SIZE),
				to_sfixed(-0.9064,1,L_SIZE),
				to_sfixed(-0.9063,1,L_SIZE),
				to_sfixed(-0.9063,1,L_SIZE),
				to_sfixed(-0.9062,1,L_SIZE),
				to_sfixed(-0.9061,1,L_SIZE),
				to_sfixed(-0.9061,1,L_SIZE),
				to_sfixed(-0.9060,1,L_SIZE),
				to_sfixed(-0.9059,1,L_SIZE),
				to_sfixed(-0.9059,1,L_SIZE),
				to_sfixed(-0.9058,1,L_SIZE),
				to_sfixed(-0.9057,1,L_SIZE),
				to_sfixed(-0.9057,1,L_SIZE),
				to_sfixed(-0.9056,1,L_SIZE),
				to_sfixed(-0.9055,1,L_SIZE),
				to_sfixed(-0.9055,1,L_SIZE),
				to_sfixed(-0.9054,1,L_SIZE),
				to_sfixed(-0.9053,1,L_SIZE),
				to_sfixed(-0.9053,1,L_SIZE),
				to_sfixed(-0.9052,1,L_SIZE),
				to_sfixed(-0.9051,1,L_SIZE),
				to_sfixed(-0.9051,1,L_SIZE),
				to_sfixed(-0.9050,1,L_SIZE),
				to_sfixed(-0.9049,1,L_SIZE),
				to_sfixed(-0.9049,1,L_SIZE),
				to_sfixed(-0.9048,1,L_SIZE),
				to_sfixed(-0.9048,1,L_SIZE),
				to_sfixed(-0.9047,1,L_SIZE),
				to_sfixed(-0.9046,1,L_SIZE),
				to_sfixed(-0.9046,1,L_SIZE),
				to_sfixed(-0.9045,1,L_SIZE),
				to_sfixed(-0.9044,1,L_SIZE),
				to_sfixed(-0.9044,1,L_SIZE),
				to_sfixed(-0.9043,1,L_SIZE),
				to_sfixed(-0.9042,1,L_SIZE),
				to_sfixed(-0.9042,1,L_SIZE),
				to_sfixed(-0.9041,1,L_SIZE),
				to_sfixed(-0.9040,1,L_SIZE),
				to_sfixed(-0.9039,1,L_SIZE),
				to_sfixed(-0.9039,1,L_SIZE),
				to_sfixed(-0.9038,1,L_SIZE),
				to_sfixed(-0.9037,1,L_SIZE),
				to_sfixed(-0.9037,1,L_SIZE),
				to_sfixed(-0.9036,1,L_SIZE),
				to_sfixed(-0.9035,1,L_SIZE),
				to_sfixed(-0.9035,1,L_SIZE),
				to_sfixed(-0.9034,1,L_SIZE),
				to_sfixed(-0.9033,1,L_SIZE),
				to_sfixed(-0.9033,1,L_SIZE),
				to_sfixed(-0.9032,1,L_SIZE),
				to_sfixed(-0.9031,1,L_SIZE),
				to_sfixed(-0.9031,1,L_SIZE),
				to_sfixed(-0.9030,1,L_SIZE),
				to_sfixed(-0.9029,1,L_SIZE),
				to_sfixed(-0.9029,1,L_SIZE),
				to_sfixed(-0.9028,1,L_SIZE),
				to_sfixed(-0.9027,1,L_SIZE),
				to_sfixed(-0.9027,1,L_SIZE),
				to_sfixed(-0.9026,1,L_SIZE),
				to_sfixed(-0.9025,1,L_SIZE),
				to_sfixed(-0.9025,1,L_SIZE),
				to_sfixed(-0.9024,1,L_SIZE),
				to_sfixed(-0.9023,1,L_SIZE),
				to_sfixed(-0.9023,1,L_SIZE),
				to_sfixed(-0.9022,1,L_SIZE),
				to_sfixed(-0.9021,1,L_SIZE),
				to_sfixed(-0.9021,1,L_SIZE),
				to_sfixed(-0.9020,1,L_SIZE),
				to_sfixed(-0.9019,1,L_SIZE),
				to_sfixed(-0.9019,1,L_SIZE),
				to_sfixed(-0.9018,1,L_SIZE),
				to_sfixed(-0.9017,1,L_SIZE),
				to_sfixed(-0.9016,1,L_SIZE),
				to_sfixed(-0.9016,1,L_SIZE),
				to_sfixed(-0.9015,1,L_SIZE),
				to_sfixed(-0.9014,1,L_SIZE),
				to_sfixed(-0.9014,1,L_SIZE),
				to_sfixed(-0.9013,1,L_SIZE),
				to_sfixed(-0.9012,1,L_SIZE),
				to_sfixed(-0.9012,1,L_SIZE),
				to_sfixed(-0.9011,1,L_SIZE),
				to_sfixed(-0.9010,1,L_SIZE),
				to_sfixed(-0.9010,1,L_SIZE),
				to_sfixed(-0.9009,1,L_SIZE),
				to_sfixed(-0.9008,1,L_SIZE),
				to_sfixed(-0.9008,1,L_SIZE),
				to_sfixed(-0.9007,1,L_SIZE),
				to_sfixed(-0.9006,1,L_SIZE),
				to_sfixed(-0.9005,1,L_SIZE),
				to_sfixed(-0.9005,1,L_SIZE),
				to_sfixed(-0.9004,1,L_SIZE),
				to_sfixed(-0.9003,1,L_SIZE),
				to_sfixed(-0.9003,1,L_SIZE),
				to_sfixed(-0.9002,1,L_SIZE),
				to_sfixed(-0.9001,1,L_SIZE),
				to_sfixed(-0.9001,1,L_SIZE),
				to_sfixed(-0.9000,1,L_SIZE),
				to_sfixed(-0.8999,1,L_SIZE),
				to_sfixed(-0.8999,1,L_SIZE),
				to_sfixed(-0.8998,1,L_SIZE),
				to_sfixed(-0.8997,1,L_SIZE),
				to_sfixed(-0.8996,1,L_SIZE),
				to_sfixed(-0.8996,1,L_SIZE),
				to_sfixed(-0.8995,1,L_SIZE),
				to_sfixed(-0.8994,1,L_SIZE),
				to_sfixed(-0.8994,1,L_SIZE),
				to_sfixed(-0.8993,1,L_SIZE),
				to_sfixed(-0.8992,1,L_SIZE),
				to_sfixed(-0.8992,1,L_SIZE),
				to_sfixed(-0.8991,1,L_SIZE),
				to_sfixed(-0.8990,1,L_SIZE),
				to_sfixed(-0.8989,1,L_SIZE),
				to_sfixed(-0.8989,1,L_SIZE),
				to_sfixed(-0.8988,1,L_SIZE),
				to_sfixed(-0.8987,1,L_SIZE),
				to_sfixed(-0.8987,1,L_SIZE),
				to_sfixed(-0.8986,1,L_SIZE),
				to_sfixed(-0.8985,1,L_SIZE),
				to_sfixed(-0.8984,1,L_SIZE),
				to_sfixed(-0.8984,1,L_SIZE),
				to_sfixed(-0.8983,1,L_SIZE),
				to_sfixed(-0.8982,1,L_SIZE),
				to_sfixed(-0.8982,1,L_SIZE),
				to_sfixed(-0.8981,1,L_SIZE),
				to_sfixed(-0.8980,1,L_SIZE),
				to_sfixed(-0.8980,1,L_SIZE),
				to_sfixed(-0.8979,1,L_SIZE),
				to_sfixed(-0.8978,1,L_SIZE),
				to_sfixed(-0.8977,1,L_SIZE),
				to_sfixed(-0.8977,1,L_SIZE),
				to_sfixed(-0.8976,1,L_SIZE),
				to_sfixed(-0.8975,1,L_SIZE),
				to_sfixed(-0.8975,1,L_SIZE),
				to_sfixed(-0.8974,1,L_SIZE),
				to_sfixed(-0.8973,1,L_SIZE),
				to_sfixed(-0.8972,1,L_SIZE),
				to_sfixed(-0.8972,1,L_SIZE),
				to_sfixed(-0.8971,1,L_SIZE),
				to_sfixed(-0.8970,1,L_SIZE),
				to_sfixed(-0.8970,1,L_SIZE),
				to_sfixed(-0.8969,1,L_SIZE),
				to_sfixed(-0.8968,1,L_SIZE),
				to_sfixed(-0.8967,1,L_SIZE),
				to_sfixed(-0.8967,1,L_SIZE),
				to_sfixed(-0.8966,1,L_SIZE),
				to_sfixed(-0.8965,1,L_SIZE),
				to_sfixed(-0.8965,1,L_SIZE),
				to_sfixed(-0.8964,1,L_SIZE),
				to_sfixed(-0.8963,1,L_SIZE),
				to_sfixed(-0.8962,1,L_SIZE),
				to_sfixed(-0.8962,1,L_SIZE),
				to_sfixed(-0.8961,1,L_SIZE),
				to_sfixed(-0.8960,1,L_SIZE),
				to_sfixed(-0.8959,1,L_SIZE),
				to_sfixed(-0.8959,1,L_SIZE),
				to_sfixed(-0.8958,1,L_SIZE),
				to_sfixed(-0.8957,1,L_SIZE),
				to_sfixed(-0.8957,1,L_SIZE),
				to_sfixed(-0.8956,1,L_SIZE),
				to_sfixed(-0.8955,1,L_SIZE),
				to_sfixed(-0.8954,1,L_SIZE),
				to_sfixed(-0.8954,1,L_SIZE),
				to_sfixed(-0.8953,1,L_SIZE),
				to_sfixed(-0.8952,1,L_SIZE),
				to_sfixed(-0.8952,1,L_SIZE),
				to_sfixed(-0.8951,1,L_SIZE),
				to_sfixed(-0.8950,1,L_SIZE),
				to_sfixed(-0.8949,1,L_SIZE),
				to_sfixed(-0.8949,1,L_SIZE),
				to_sfixed(-0.8948,1,L_SIZE),
				to_sfixed(-0.8947,1,L_SIZE),
				to_sfixed(-0.8946,1,L_SIZE),
				to_sfixed(-0.8946,1,L_SIZE),
				to_sfixed(-0.8945,1,L_SIZE),
				to_sfixed(-0.8944,1,L_SIZE),
				to_sfixed(-0.8943,1,L_SIZE),
				to_sfixed(-0.8943,1,L_SIZE),
				to_sfixed(-0.8942,1,L_SIZE),
				to_sfixed(-0.8941,1,L_SIZE),
				to_sfixed(-0.8941,1,L_SIZE),
				to_sfixed(-0.8940,1,L_SIZE),
				to_sfixed(-0.8939,1,L_SIZE),
				to_sfixed(-0.8938,1,L_SIZE),
				to_sfixed(-0.8938,1,L_SIZE),
				to_sfixed(-0.8937,1,L_SIZE),
				to_sfixed(-0.8936,1,L_SIZE),
				to_sfixed(-0.8935,1,L_SIZE),
				to_sfixed(-0.8935,1,L_SIZE),
				to_sfixed(-0.8934,1,L_SIZE),
				to_sfixed(-0.8933,1,L_SIZE),
				to_sfixed(-0.8932,1,L_SIZE),
				to_sfixed(-0.8932,1,L_SIZE),
				to_sfixed(-0.8931,1,L_SIZE),
				to_sfixed(-0.8930,1,L_SIZE),
				to_sfixed(-0.8929,1,L_SIZE),
				to_sfixed(-0.8929,1,L_SIZE),
				to_sfixed(-0.8928,1,L_SIZE),
				to_sfixed(-0.8927,1,L_SIZE),
				to_sfixed(-0.8926,1,L_SIZE),
				to_sfixed(-0.8926,1,L_SIZE),
				to_sfixed(-0.8925,1,L_SIZE),
				to_sfixed(-0.8924,1,L_SIZE),
				to_sfixed(-0.8924,1,L_SIZE),
				to_sfixed(-0.8923,1,L_SIZE),
				to_sfixed(-0.8922,1,L_SIZE),
				to_sfixed(-0.8921,1,L_SIZE),
				to_sfixed(-0.8921,1,L_SIZE),
				to_sfixed(-0.8920,1,L_SIZE),
				to_sfixed(-0.8919,1,L_SIZE),
				to_sfixed(-0.8918,1,L_SIZE),
				to_sfixed(-0.8918,1,L_SIZE),
				to_sfixed(-0.8917,1,L_SIZE),
				to_sfixed(-0.8916,1,L_SIZE),
				to_sfixed(-0.8915,1,L_SIZE),
				to_sfixed(-0.8915,1,L_SIZE),
				to_sfixed(-0.8914,1,L_SIZE),
				to_sfixed(-0.8913,1,L_SIZE),
				to_sfixed(-0.8912,1,L_SIZE),
				to_sfixed(-0.8912,1,L_SIZE),
				to_sfixed(-0.8911,1,L_SIZE),
				to_sfixed(-0.8910,1,L_SIZE),
				to_sfixed(-0.8909,1,L_SIZE),
				to_sfixed(-0.8908,1,L_SIZE),
				to_sfixed(-0.8908,1,L_SIZE),
				to_sfixed(-0.8907,1,L_SIZE),
				to_sfixed(-0.8906,1,L_SIZE),
				to_sfixed(-0.8905,1,L_SIZE),
				to_sfixed(-0.8905,1,L_SIZE),
				to_sfixed(-0.8904,1,L_SIZE),
				to_sfixed(-0.8903,1,L_SIZE),
				to_sfixed(-0.8902,1,L_SIZE),
				to_sfixed(-0.8902,1,L_SIZE),
				to_sfixed(-0.8901,1,L_SIZE),
				to_sfixed(-0.8900,1,L_SIZE),
				to_sfixed(-0.8899,1,L_SIZE),
				to_sfixed(-0.8899,1,L_SIZE),
				to_sfixed(-0.8898,1,L_SIZE),
				to_sfixed(-0.8897,1,L_SIZE),
				to_sfixed(-0.8896,1,L_SIZE),
				to_sfixed(-0.8896,1,L_SIZE),
				to_sfixed(-0.8895,1,L_SIZE),
				to_sfixed(-0.8894,1,L_SIZE),
				to_sfixed(-0.8893,1,L_SIZE),
				to_sfixed(-0.8893,1,L_SIZE),
				to_sfixed(-0.8892,1,L_SIZE),
				to_sfixed(-0.8891,1,L_SIZE),
				to_sfixed(-0.8890,1,L_SIZE),
				to_sfixed(-0.8889,1,L_SIZE),
				to_sfixed(-0.8889,1,L_SIZE),
				to_sfixed(-0.8888,1,L_SIZE),
				to_sfixed(-0.8887,1,L_SIZE),
				to_sfixed(-0.8886,1,L_SIZE),
				to_sfixed(-0.8886,1,L_SIZE),
				to_sfixed(-0.8885,1,L_SIZE),
				to_sfixed(-0.8884,1,L_SIZE),
				to_sfixed(-0.8883,1,L_SIZE),
				to_sfixed(-0.8883,1,L_SIZE),
				to_sfixed(-0.8882,1,L_SIZE),
				to_sfixed(-0.8881,1,L_SIZE),
				to_sfixed(-0.8880,1,L_SIZE),
				to_sfixed(-0.8879,1,L_SIZE),
				to_sfixed(-0.8879,1,L_SIZE),
				to_sfixed(-0.8878,1,L_SIZE),
				to_sfixed(-0.8877,1,L_SIZE),
				to_sfixed(-0.8876,1,L_SIZE),
				to_sfixed(-0.8876,1,L_SIZE),
				to_sfixed(-0.8875,1,L_SIZE),
				to_sfixed(-0.8874,1,L_SIZE),
				to_sfixed(-0.8873,1,L_SIZE),
				to_sfixed(-0.8872,1,L_SIZE),
				to_sfixed(-0.8872,1,L_SIZE),
				to_sfixed(-0.8871,1,L_SIZE),
				to_sfixed(-0.8870,1,L_SIZE),
				to_sfixed(-0.8869,1,L_SIZE),
				to_sfixed(-0.8869,1,L_SIZE),
				to_sfixed(-0.8868,1,L_SIZE),
				to_sfixed(-0.8867,1,L_SIZE),
				to_sfixed(-0.8866,1,L_SIZE),
				to_sfixed(-0.8865,1,L_SIZE),
				to_sfixed(-0.8865,1,L_SIZE),
				to_sfixed(-0.8864,1,L_SIZE),
				to_sfixed(-0.8863,1,L_SIZE),
				to_sfixed(-0.8862,1,L_SIZE),
				to_sfixed(-0.8861,1,L_SIZE),
				to_sfixed(-0.8861,1,L_SIZE),
				to_sfixed(-0.8860,1,L_SIZE),
				to_sfixed(-0.8859,1,L_SIZE),
				to_sfixed(-0.8858,1,L_SIZE),
				to_sfixed(-0.8858,1,L_SIZE),
				to_sfixed(-0.8857,1,L_SIZE),
				to_sfixed(-0.8856,1,L_SIZE),
				to_sfixed(-0.8855,1,L_SIZE),
				to_sfixed(-0.8854,1,L_SIZE),
				to_sfixed(-0.8854,1,L_SIZE),
				to_sfixed(-0.8853,1,L_SIZE),
				to_sfixed(-0.8852,1,L_SIZE),
				to_sfixed(-0.8851,1,L_SIZE),
				to_sfixed(-0.8850,1,L_SIZE),
				to_sfixed(-0.8850,1,L_SIZE),
				to_sfixed(-0.8849,1,L_SIZE),
				to_sfixed(-0.8848,1,L_SIZE),
				to_sfixed(-0.8847,1,L_SIZE),
				to_sfixed(-0.8846,1,L_SIZE),
				to_sfixed(-0.8846,1,L_SIZE),
				to_sfixed(-0.8845,1,L_SIZE),
				to_sfixed(-0.8844,1,L_SIZE),
				to_sfixed(-0.8843,1,L_SIZE),
				to_sfixed(-0.8842,1,L_SIZE),
				to_sfixed(-0.8842,1,L_SIZE),
				to_sfixed(-0.8841,1,L_SIZE),
				to_sfixed(-0.8840,1,L_SIZE),
				to_sfixed(-0.8839,1,L_SIZE),
				to_sfixed(-0.8838,1,L_SIZE),
				to_sfixed(-0.8838,1,L_SIZE),
				to_sfixed(-0.8837,1,L_SIZE),
				to_sfixed(-0.8836,1,L_SIZE),
				to_sfixed(-0.8835,1,L_SIZE),
				to_sfixed(-0.8834,1,L_SIZE),
				to_sfixed(-0.8834,1,L_SIZE),
				to_sfixed(-0.8833,1,L_SIZE),
				to_sfixed(-0.8832,1,L_SIZE),
				to_sfixed(-0.8831,1,L_SIZE),
				to_sfixed(-0.8830,1,L_SIZE),
				to_sfixed(-0.8830,1,L_SIZE),
				to_sfixed(-0.8829,1,L_SIZE),
				to_sfixed(-0.8828,1,L_SIZE),
				to_sfixed(-0.8827,1,L_SIZE),
				to_sfixed(-0.8826,1,L_SIZE),
				to_sfixed(-0.8826,1,L_SIZE),
				to_sfixed(-0.8825,1,L_SIZE),
				to_sfixed(-0.8824,1,L_SIZE),
				to_sfixed(-0.8823,1,L_SIZE),
				to_sfixed(-0.8822,1,L_SIZE),
				to_sfixed(-0.8821,1,L_SIZE),
				to_sfixed(-0.8821,1,L_SIZE),
				to_sfixed(-0.8820,1,L_SIZE),
				to_sfixed(-0.8819,1,L_SIZE),
				to_sfixed(-0.8818,1,L_SIZE),
				to_sfixed(-0.8817,1,L_SIZE),
				to_sfixed(-0.8817,1,L_SIZE),
				to_sfixed(-0.8816,1,L_SIZE),
				to_sfixed(-0.8815,1,L_SIZE),
				to_sfixed(-0.8814,1,L_SIZE),
				to_sfixed(-0.8813,1,L_SIZE),
				to_sfixed(-0.8813,1,L_SIZE),
				to_sfixed(-0.8812,1,L_SIZE),
				to_sfixed(-0.8811,1,L_SIZE),
				to_sfixed(-0.8810,1,L_SIZE),
				to_sfixed(-0.8809,1,L_SIZE),
				to_sfixed(-0.8808,1,L_SIZE),
				to_sfixed(-0.8808,1,L_SIZE),
				to_sfixed(-0.8807,1,L_SIZE),
				to_sfixed(-0.8806,1,L_SIZE),
				to_sfixed(-0.8805,1,L_SIZE),
				to_sfixed(-0.8804,1,L_SIZE),
				to_sfixed(-0.8803,1,L_SIZE),
				to_sfixed(-0.8803,1,L_SIZE),
				to_sfixed(-0.8802,1,L_SIZE),
				to_sfixed(-0.8801,1,L_SIZE),
				to_sfixed(-0.8800,1,L_SIZE),
				to_sfixed(-0.8799,1,L_SIZE),
				to_sfixed(-0.8799,1,L_SIZE),
				to_sfixed(-0.8798,1,L_SIZE),
				to_sfixed(-0.8797,1,L_SIZE),
				to_sfixed(-0.8796,1,L_SIZE),
				to_sfixed(-0.8795,1,L_SIZE),
				to_sfixed(-0.8794,1,L_SIZE),
				to_sfixed(-0.8794,1,L_SIZE),
				to_sfixed(-0.8793,1,L_SIZE),
				to_sfixed(-0.8792,1,L_SIZE),
				to_sfixed(-0.8791,1,L_SIZE),
				to_sfixed(-0.8790,1,L_SIZE),
				to_sfixed(-0.8789,1,L_SIZE),
				to_sfixed(-0.8789,1,L_SIZE),
				to_sfixed(-0.8788,1,L_SIZE),
				to_sfixed(-0.8787,1,L_SIZE),
				to_sfixed(-0.8786,1,L_SIZE),
				to_sfixed(-0.8785,1,L_SIZE),
				to_sfixed(-0.8784,1,L_SIZE),
				to_sfixed(-0.8784,1,L_SIZE),
				to_sfixed(-0.8783,1,L_SIZE),
				to_sfixed(-0.8782,1,L_SIZE),
				to_sfixed(-0.8781,1,L_SIZE),
				to_sfixed(-0.8780,1,L_SIZE),
				to_sfixed(-0.8779,1,L_SIZE),
				to_sfixed(-0.8779,1,L_SIZE),
				to_sfixed(-0.8778,1,L_SIZE),
				to_sfixed(-0.8777,1,L_SIZE),
				to_sfixed(-0.8776,1,L_SIZE),
				to_sfixed(-0.8775,1,L_SIZE),
				to_sfixed(-0.8774,1,L_SIZE),
				to_sfixed(-0.8773,1,L_SIZE),
				to_sfixed(-0.8773,1,L_SIZE),
				to_sfixed(-0.8772,1,L_SIZE),
				to_sfixed(-0.8771,1,L_SIZE),
				to_sfixed(-0.8770,1,L_SIZE),
				to_sfixed(-0.8769,1,L_SIZE),
				to_sfixed(-0.8768,1,L_SIZE),
				to_sfixed(-0.8768,1,L_SIZE),
				to_sfixed(-0.8767,1,L_SIZE),
				to_sfixed(-0.8766,1,L_SIZE),
				to_sfixed(-0.8765,1,L_SIZE),
				to_sfixed(-0.8764,1,L_SIZE),
				to_sfixed(-0.8763,1,L_SIZE),
				to_sfixed(-0.8762,1,L_SIZE),
				to_sfixed(-0.8762,1,L_SIZE),
				to_sfixed(-0.8761,1,L_SIZE),
				to_sfixed(-0.8760,1,L_SIZE),
				to_sfixed(-0.8759,1,L_SIZE),
				to_sfixed(-0.8758,1,L_SIZE),
				to_sfixed(-0.8757,1,L_SIZE),
				to_sfixed(-0.8757,1,L_SIZE),
				to_sfixed(-0.8756,1,L_SIZE),
				to_sfixed(-0.8755,1,L_SIZE),
				to_sfixed(-0.8754,1,L_SIZE),
				to_sfixed(-0.8753,1,L_SIZE),
				to_sfixed(-0.8752,1,L_SIZE),
				to_sfixed(-0.8751,1,L_SIZE),
				to_sfixed(-0.8751,1,L_SIZE),
				to_sfixed(-0.8750,1,L_SIZE),
				to_sfixed(-0.8749,1,L_SIZE),
				to_sfixed(-0.8748,1,L_SIZE),
				to_sfixed(-0.8747,1,L_SIZE),
				to_sfixed(-0.8746,1,L_SIZE),
				to_sfixed(-0.8745,1,L_SIZE),
				to_sfixed(-0.8745,1,L_SIZE),
				to_sfixed(-0.8744,1,L_SIZE),
				to_sfixed(-0.8743,1,L_SIZE),
				to_sfixed(-0.8742,1,L_SIZE),
				to_sfixed(-0.8741,1,L_SIZE),
				to_sfixed(-0.8740,1,L_SIZE),
				to_sfixed(-0.8739,1,L_SIZE),
				to_sfixed(-0.8738,1,L_SIZE),
				to_sfixed(-0.8738,1,L_SIZE),
				to_sfixed(-0.8737,1,L_SIZE),
				to_sfixed(-0.8736,1,L_SIZE),
				to_sfixed(-0.8735,1,L_SIZE),
				to_sfixed(-0.8734,1,L_SIZE),
				to_sfixed(-0.8733,1,L_SIZE),
				to_sfixed(-0.8732,1,L_SIZE),
				to_sfixed(-0.8732,1,L_SIZE),
				to_sfixed(-0.8731,1,L_SIZE),
				to_sfixed(-0.8730,1,L_SIZE),
				to_sfixed(-0.8729,1,L_SIZE),
				to_sfixed(-0.8728,1,L_SIZE),
				to_sfixed(-0.8727,1,L_SIZE),
				to_sfixed(-0.8726,1,L_SIZE),
				to_sfixed(-0.8725,1,L_SIZE),
				to_sfixed(-0.8725,1,L_SIZE),
				to_sfixed(-0.8724,1,L_SIZE),
				to_sfixed(-0.8723,1,L_SIZE),
				to_sfixed(-0.8722,1,L_SIZE),
				to_sfixed(-0.8721,1,L_SIZE),
				to_sfixed(-0.8720,1,L_SIZE),
				to_sfixed(-0.8719,1,L_SIZE),
				to_sfixed(-0.8718,1,L_SIZE),
				to_sfixed(-0.8718,1,L_SIZE),
				to_sfixed(-0.8717,1,L_SIZE),
				to_sfixed(-0.8716,1,L_SIZE),
				to_sfixed(-0.8715,1,L_SIZE),
				to_sfixed(-0.8714,1,L_SIZE),
				to_sfixed(-0.8713,1,L_SIZE),
				to_sfixed(-0.8712,1,L_SIZE),
				to_sfixed(-0.8711,1,L_SIZE),
				to_sfixed(-0.8710,1,L_SIZE),
				to_sfixed(-0.8710,1,L_SIZE),
				to_sfixed(-0.8709,1,L_SIZE),
				to_sfixed(-0.8708,1,L_SIZE),
				to_sfixed(-0.8707,1,L_SIZE),
				to_sfixed(-0.8706,1,L_SIZE),
				to_sfixed(-0.8705,1,L_SIZE),
				to_sfixed(-0.8704,1,L_SIZE),
				to_sfixed(-0.8703,1,L_SIZE),
				to_sfixed(-0.8702,1,L_SIZE),
				to_sfixed(-0.8702,1,L_SIZE),
				to_sfixed(-0.8701,1,L_SIZE),
				to_sfixed(-0.8700,1,L_SIZE),
				to_sfixed(-0.8699,1,L_SIZE),
				to_sfixed(-0.8698,1,L_SIZE),
				to_sfixed(-0.8697,1,L_SIZE),
				to_sfixed(-0.8696,1,L_SIZE),
				to_sfixed(-0.8695,1,L_SIZE),
				to_sfixed(-0.8694,1,L_SIZE),
				to_sfixed(-0.8694,1,L_SIZE),
				to_sfixed(-0.8693,1,L_SIZE),
				to_sfixed(-0.8692,1,L_SIZE),
				to_sfixed(-0.8691,1,L_SIZE),
				to_sfixed(-0.8690,1,L_SIZE),
				to_sfixed(-0.8689,1,L_SIZE),
				to_sfixed(-0.8688,1,L_SIZE),
				to_sfixed(-0.8687,1,L_SIZE),
				to_sfixed(-0.8686,1,L_SIZE),
				to_sfixed(-0.8686,1,L_SIZE),
				to_sfixed(-0.8685,1,L_SIZE),
				to_sfixed(-0.8684,1,L_SIZE),
				to_sfixed(-0.8683,1,L_SIZE),
				to_sfixed(-0.8682,1,L_SIZE),
				to_sfixed(-0.8681,1,L_SIZE),
				to_sfixed(-0.8680,1,L_SIZE),
				to_sfixed(-0.8679,1,L_SIZE),
				to_sfixed(-0.8678,1,L_SIZE),
				to_sfixed(-0.8677,1,L_SIZE),
				to_sfixed(-0.8676,1,L_SIZE),
				to_sfixed(-0.8676,1,L_SIZE),
				to_sfixed(-0.8675,1,L_SIZE),
				to_sfixed(-0.8674,1,L_SIZE),
				to_sfixed(-0.8673,1,L_SIZE),
				to_sfixed(-0.8672,1,L_SIZE),
				to_sfixed(-0.8671,1,L_SIZE),
				to_sfixed(-0.8670,1,L_SIZE),
				to_sfixed(-0.8669,1,L_SIZE),
				to_sfixed(-0.8668,1,L_SIZE),
				to_sfixed(-0.8667,1,L_SIZE),
				to_sfixed(-0.8666,1,L_SIZE),
				to_sfixed(-0.8666,1,L_SIZE),
				to_sfixed(-0.8665,1,L_SIZE),
				to_sfixed(-0.8664,1,L_SIZE),
				to_sfixed(-0.8663,1,L_SIZE),
				to_sfixed(-0.8662,1,L_SIZE),
				to_sfixed(-0.8661,1,L_SIZE),
				to_sfixed(-0.8660,1,L_SIZE),
				to_sfixed(-0.8659,1,L_SIZE),
				to_sfixed(-0.8658,1,L_SIZE),
				to_sfixed(-0.8657,1,L_SIZE),
				to_sfixed(-0.8656,1,L_SIZE),
				to_sfixed(-0.8656,1,L_SIZE),
				to_sfixed(-0.8655,1,L_SIZE),
				to_sfixed(-0.8654,1,L_SIZE),
				to_sfixed(-0.8653,1,L_SIZE),
				to_sfixed(-0.8652,1,L_SIZE),
				to_sfixed(-0.8651,1,L_SIZE),
				to_sfixed(-0.8650,1,L_SIZE),
				to_sfixed(-0.8649,1,L_SIZE),
				to_sfixed(-0.8648,1,L_SIZE),
				to_sfixed(-0.8647,1,L_SIZE),
				to_sfixed(-0.8646,1,L_SIZE),
				to_sfixed(-0.8645,1,L_SIZE),
				to_sfixed(-0.8644,1,L_SIZE),
				to_sfixed(-0.8644,1,L_SIZE),
				to_sfixed(-0.8643,1,L_SIZE),
				to_sfixed(-0.8642,1,L_SIZE),
				to_sfixed(-0.8641,1,L_SIZE),
				to_sfixed(-0.8640,1,L_SIZE),
				to_sfixed(-0.8639,1,L_SIZE),
				to_sfixed(-0.8638,1,L_SIZE),
				to_sfixed(-0.8637,1,L_SIZE),
				to_sfixed(-0.8636,1,L_SIZE),
				to_sfixed(-0.8635,1,L_SIZE),
				to_sfixed(-0.8634,1,L_SIZE),
				to_sfixed(-0.8633,1,L_SIZE),
				to_sfixed(-0.8632,1,L_SIZE),
				to_sfixed(-0.8631,1,L_SIZE),
				to_sfixed(-0.8630,1,L_SIZE),
				to_sfixed(-0.8630,1,L_SIZE),
				to_sfixed(-0.8629,1,L_SIZE),
				to_sfixed(-0.8628,1,L_SIZE),
				to_sfixed(-0.8627,1,L_SIZE),
				to_sfixed(-0.8626,1,L_SIZE),
				to_sfixed(-0.8625,1,L_SIZE),
				to_sfixed(-0.8624,1,L_SIZE),
				to_sfixed(-0.8623,1,L_SIZE),
				to_sfixed(-0.8622,1,L_SIZE),
				to_sfixed(-0.8621,1,L_SIZE),
				to_sfixed(-0.8620,1,L_SIZE),
				to_sfixed(-0.8619,1,L_SIZE),
				to_sfixed(-0.8618,1,L_SIZE),
				to_sfixed(-0.8617,1,L_SIZE),
				to_sfixed(-0.8616,1,L_SIZE),
				to_sfixed(-0.8615,1,L_SIZE),
				to_sfixed(-0.8615,1,L_SIZE),
				to_sfixed(-0.8614,1,L_SIZE),
				to_sfixed(-0.8613,1,L_SIZE),
				to_sfixed(-0.8612,1,L_SIZE),
				to_sfixed(-0.8611,1,L_SIZE),
				to_sfixed(-0.8610,1,L_SIZE),
				to_sfixed(-0.8609,1,L_SIZE),
				to_sfixed(-0.8608,1,L_SIZE),
				to_sfixed(-0.8607,1,L_SIZE),
				to_sfixed(-0.8606,1,L_SIZE),
				to_sfixed(-0.8605,1,L_SIZE),
				to_sfixed(-0.8604,1,L_SIZE),
				to_sfixed(-0.8603,1,L_SIZE),
				to_sfixed(-0.8602,1,L_SIZE),
				to_sfixed(-0.8601,1,L_SIZE),
				to_sfixed(-0.8600,1,L_SIZE),
				to_sfixed(-0.8599,1,L_SIZE),
				to_sfixed(-0.8598,1,L_SIZE),
				to_sfixed(-0.8597,1,L_SIZE),
				to_sfixed(-0.8596,1,L_SIZE),
				to_sfixed(-0.8596,1,L_SIZE),
				to_sfixed(-0.8595,1,L_SIZE),
				to_sfixed(-0.8594,1,L_SIZE),
				to_sfixed(-0.8593,1,L_SIZE),
				to_sfixed(-0.8592,1,L_SIZE),
				to_sfixed(-0.8591,1,L_SIZE),
				to_sfixed(-0.8590,1,L_SIZE),
				to_sfixed(-0.8589,1,L_SIZE),
				to_sfixed(-0.8588,1,L_SIZE),
				to_sfixed(-0.8587,1,L_SIZE),
				to_sfixed(-0.8586,1,L_SIZE),
				to_sfixed(-0.8585,1,L_SIZE),
				to_sfixed(-0.8584,1,L_SIZE),
				to_sfixed(-0.8583,1,L_SIZE),
				to_sfixed(-0.8582,1,L_SIZE),
				to_sfixed(-0.8581,1,L_SIZE),
				to_sfixed(-0.8580,1,L_SIZE),
				to_sfixed(-0.8579,1,L_SIZE),
				to_sfixed(-0.8578,1,L_SIZE),
				to_sfixed(-0.8577,1,L_SIZE),
				to_sfixed(-0.8576,1,L_SIZE),
				to_sfixed(-0.8575,1,L_SIZE),
				to_sfixed(-0.8574,1,L_SIZE),
				to_sfixed(-0.8573,1,L_SIZE),
				to_sfixed(-0.8572,1,L_SIZE),
				to_sfixed(-0.8571,1,L_SIZE),
				to_sfixed(-0.8570,1,L_SIZE),
				to_sfixed(-0.8569,1,L_SIZE),
				to_sfixed(-0.8569,1,L_SIZE),
				to_sfixed(-0.8568,1,L_SIZE),
				to_sfixed(-0.8567,1,L_SIZE),
				to_sfixed(-0.8566,1,L_SIZE),
				to_sfixed(-0.8565,1,L_SIZE),
				to_sfixed(-0.8564,1,L_SIZE),
				to_sfixed(-0.8563,1,L_SIZE),
				to_sfixed(-0.8562,1,L_SIZE),
				to_sfixed(-0.8561,1,L_SIZE),
				to_sfixed(-0.8560,1,L_SIZE),
				to_sfixed(-0.8559,1,L_SIZE),
				to_sfixed(-0.8558,1,L_SIZE),
				to_sfixed(-0.8557,1,L_SIZE),
				to_sfixed(-0.8556,1,L_SIZE),
				to_sfixed(-0.8555,1,L_SIZE),
				to_sfixed(-0.8554,1,L_SIZE),
				to_sfixed(-0.8553,1,L_SIZE),
				to_sfixed(-0.8552,1,L_SIZE),
				to_sfixed(-0.8551,1,L_SIZE),
				to_sfixed(-0.8550,1,L_SIZE),
				to_sfixed(-0.8549,1,L_SIZE),
				to_sfixed(-0.8548,1,L_SIZE),
				to_sfixed(-0.8547,1,L_SIZE),
				to_sfixed(-0.8546,1,L_SIZE),
				to_sfixed(-0.8545,1,L_SIZE),
				to_sfixed(-0.8544,1,L_SIZE),
				to_sfixed(-0.8543,1,L_SIZE),
				to_sfixed(-0.8542,1,L_SIZE),
				to_sfixed(-0.8541,1,L_SIZE),
				to_sfixed(-0.8540,1,L_SIZE),
				to_sfixed(-0.8539,1,L_SIZE),
				to_sfixed(-0.8538,1,L_SIZE),
				to_sfixed(-0.8537,1,L_SIZE),
				to_sfixed(-0.8536,1,L_SIZE),
				to_sfixed(-0.8535,1,L_SIZE),
				to_sfixed(-0.8534,1,L_SIZE),
				to_sfixed(-0.8533,1,L_SIZE),
				to_sfixed(-0.8532,1,L_SIZE),
				to_sfixed(-0.8531,1,L_SIZE),
				to_sfixed(-0.8530,1,L_SIZE),
				to_sfixed(-0.8529,1,L_SIZE),
				to_sfixed(-0.8528,1,L_SIZE),
				to_sfixed(-0.8527,1,L_SIZE),
				to_sfixed(-0.8526,1,L_SIZE),
				to_sfixed(-0.8525,1,L_SIZE),
				to_sfixed(-0.8524,1,L_SIZE),
				to_sfixed(-0.8523,1,L_SIZE),
				to_sfixed(-0.8522,1,L_SIZE),
				to_sfixed(-0.8521,1,L_SIZE),
				to_sfixed(-0.8520,1,L_SIZE),
				to_sfixed(-0.8519,1,L_SIZE),
				to_sfixed(-0.8518,1,L_SIZE),
				to_sfixed(-0.8517,1,L_SIZE),
				to_sfixed(-0.8516,1,L_SIZE),
				to_sfixed(-0.8515,1,L_SIZE),
				to_sfixed(-0.8514,1,L_SIZE),
				to_sfixed(-0.8513,1,L_SIZE),
				to_sfixed(-0.8512,1,L_SIZE),
				to_sfixed(-0.8511,1,L_SIZE),
				to_sfixed(-0.8510,1,L_SIZE),
				to_sfixed(-0.8509,1,L_SIZE),
				to_sfixed(-0.8508,1,L_SIZE),
				to_sfixed(-0.8507,1,L_SIZE),
				to_sfixed(-0.8506,1,L_SIZE),
				to_sfixed(-0.8505,1,L_SIZE),
				to_sfixed(-0.8504,1,L_SIZE),
				to_sfixed(-0.8503,1,L_SIZE),
				to_sfixed(-0.8502,1,L_SIZE),
				to_sfixed(-0.8501,1,L_SIZE),
				to_sfixed(-0.8500,1,L_SIZE),
				to_sfixed(-0.8499,1,L_SIZE),
				to_sfixed(-0.8498,1,L_SIZE),
				to_sfixed(-0.8497,1,L_SIZE),
				to_sfixed(-0.8496,1,L_SIZE),
				to_sfixed(-0.8495,1,L_SIZE),
				to_sfixed(-0.8494,1,L_SIZE),
				to_sfixed(-0.8493,1,L_SIZE),
				to_sfixed(-0.8492,1,L_SIZE),
				to_sfixed(-0.8491,1,L_SIZE),
				to_sfixed(-0.8490,1,L_SIZE),
				to_sfixed(-0.8489,1,L_SIZE),
				to_sfixed(-0.8488,1,L_SIZE),
				to_sfixed(-0.8487,1,L_SIZE),
				to_sfixed(-0.8486,1,L_SIZE),
				to_sfixed(-0.8485,1,L_SIZE),
				to_sfixed(-0.8484,1,L_SIZE),
				to_sfixed(-0.8482,1,L_SIZE),
				to_sfixed(-0.8481,1,L_SIZE),
				to_sfixed(-0.8480,1,L_SIZE),
				to_sfixed(-0.8479,1,L_SIZE),
				to_sfixed(-0.8478,1,L_SIZE),
				to_sfixed(-0.8477,1,L_SIZE),
				to_sfixed(-0.8476,1,L_SIZE),
				to_sfixed(-0.8475,1,L_SIZE),
				to_sfixed(-0.8474,1,L_SIZE),
				to_sfixed(-0.8473,1,L_SIZE),
				to_sfixed(-0.8472,1,L_SIZE),
				to_sfixed(-0.8471,1,L_SIZE),
				to_sfixed(-0.8470,1,L_SIZE),
				to_sfixed(-0.8469,1,L_SIZE),
				to_sfixed(-0.8468,1,L_SIZE),
				to_sfixed(-0.8467,1,L_SIZE),
				to_sfixed(-0.8466,1,L_SIZE),
				to_sfixed(-0.8465,1,L_SIZE),
				to_sfixed(-0.8464,1,L_SIZE),
				to_sfixed(-0.8463,1,L_SIZE),
				to_sfixed(-0.8462,1,L_SIZE),
				to_sfixed(-0.8461,1,L_SIZE),
				to_sfixed(-0.8460,1,L_SIZE),
				to_sfixed(-0.8459,1,L_SIZE),
				to_sfixed(-0.8458,1,L_SIZE),
				to_sfixed(-0.8457,1,L_SIZE),
				to_sfixed(-0.8456,1,L_SIZE),
				to_sfixed(-0.8455,1,L_SIZE),
				to_sfixed(-0.8453,1,L_SIZE),
				to_sfixed(-0.8452,1,L_SIZE),
				to_sfixed(-0.8451,1,L_SIZE),
				to_sfixed(-0.8450,1,L_SIZE),
				to_sfixed(-0.8449,1,L_SIZE),
				to_sfixed(-0.8448,1,L_SIZE),
				to_sfixed(-0.8447,1,L_SIZE),
				to_sfixed(-0.8446,1,L_SIZE),
				to_sfixed(-0.8445,1,L_SIZE),
				to_sfixed(-0.8444,1,L_SIZE),
				to_sfixed(-0.8443,1,L_SIZE),
				to_sfixed(-0.8442,1,L_SIZE),
				to_sfixed(-0.8441,1,L_SIZE),
				to_sfixed(-0.8440,1,L_SIZE),
				to_sfixed(-0.8439,1,L_SIZE),
				to_sfixed(-0.8438,1,L_SIZE),
				to_sfixed(-0.8437,1,L_SIZE),
				to_sfixed(-0.8436,1,L_SIZE),
				to_sfixed(-0.8435,1,L_SIZE),
				to_sfixed(-0.8434,1,L_SIZE),
				to_sfixed(-0.8432,1,L_SIZE),
				to_sfixed(-0.8431,1,L_SIZE),
				to_sfixed(-0.8430,1,L_SIZE),
				to_sfixed(-0.8429,1,L_SIZE),
				to_sfixed(-0.8428,1,L_SIZE),
				to_sfixed(-0.8427,1,L_SIZE),
				to_sfixed(-0.8426,1,L_SIZE),
				to_sfixed(-0.8425,1,L_SIZE),
				to_sfixed(-0.8424,1,L_SIZE),
				to_sfixed(-0.8423,1,L_SIZE),
				to_sfixed(-0.8422,1,L_SIZE),
				to_sfixed(-0.8421,1,L_SIZE),
				to_sfixed(-0.8420,1,L_SIZE),
				to_sfixed(-0.8419,1,L_SIZE),
				to_sfixed(-0.8418,1,L_SIZE),
				to_sfixed(-0.8417,1,L_SIZE),
				to_sfixed(-0.8415,1,L_SIZE),
				to_sfixed(-0.8414,1,L_SIZE),
				to_sfixed(-0.8413,1,L_SIZE),
				to_sfixed(-0.8412,1,L_SIZE),
				to_sfixed(-0.8411,1,L_SIZE),
				to_sfixed(-0.8410,1,L_SIZE),
				to_sfixed(-0.8409,1,L_SIZE),
				to_sfixed(-0.8408,1,L_SIZE),
				to_sfixed(-0.8407,1,L_SIZE),
				to_sfixed(-0.8406,1,L_SIZE),
				to_sfixed(-0.8405,1,L_SIZE),
				to_sfixed(-0.8404,1,L_SIZE),
				to_sfixed(-0.8403,1,L_SIZE),
				to_sfixed(-0.8401,1,L_SIZE),
				to_sfixed(-0.8400,1,L_SIZE),
				to_sfixed(-0.8399,1,L_SIZE),
				to_sfixed(-0.8398,1,L_SIZE),
				to_sfixed(-0.8397,1,L_SIZE),
				to_sfixed(-0.8396,1,L_SIZE),
				to_sfixed(-0.8395,1,L_SIZE),
				to_sfixed(-0.8394,1,L_SIZE),
				to_sfixed(-0.8393,1,L_SIZE),
				to_sfixed(-0.8392,1,L_SIZE),
				to_sfixed(-0.8391,1,L_SIZE),
				to_sfixed(-0.8390,1,L_SIZE),
				to_sfixed(-0.8389,1,L_SIZE),
				to_sfixed(-0.8387,1,L_SIZE),
				to_sfixed(-0.8386,1,L_SIZE),
				to_sfixed(-0.8385,1,L_SIZE),
				to_sfixed(-0.8384,1,L_SIZE),
				to_sfixed(-0.8383,1,L_SIZE),
				to_sfixed(-0.8382,1,L_SIZE),
				to_sfixed(-0.8381,1,L_SIZE),
				to_sfixed(-0.8380,1,L_SIZE),
				to_sfixed(-0.8379,1,L_SIZE),
				to_sfixed(-0.8378,1,L_SIZE),
				to_sfixed(-0.8377,1,L_SIZE),
				to_sfixed(-0.8375,1,L_SIZE),
				to_sfixed(-0.8374,1,L_SIZE),
				to_sfixed(-0.8373,1,L_SIZE),
				to_sfixed(-0.8372,1,L_SIZE),
				to_sfixed(-0.8371,1,L_SIZE),
				to_sfixed(-0.8370,1,L_SIZE),
				to_sfixed(-0.8369,1,L_SIZE),
				to_sfixed(-0.8368,1,L_SIZE),
				to_sfixed(-0.8367,1,L_SIZE),
				to_sfixed(-0.8366,1,L_SIZE),
				to_sfixed(-0.8364,1,L_SIZE),
				to_sfixed(-0.8363,1,L_SIZE),
				to_sfixed(-0.8362,1,L_SIZE),
				to_sfixed(-0.8361,1,L_SIZE),
				to_sfixed(-0.8360,1,L_SIZE),
				to_sfixed(-0.8359,1,L_SIZE),
				to_sfixed(-0.8358,1,L_SIZE),
				to_sfixed(-0.8357,1,L_SIZE),
				to_sfixed(-0.8356,1,L_SIZE),
				to_sfixed(-0.8355,1,L_SIZE),
				to_sfixed(-0.8353,1,L_SIZE),
				to_sfixed(-0.8352,1,L_SIZE),
				to_sfixed(-0.8351,1,L_SIZE),
				to_sfixed(-0.8350,1,L_SIZE),
				to_sfixed(-0.8349,1,L_SIZE),
				to_sfixed(-0.8348,1,L_SIZE),
				to_sfixed(-0.8347,1,L_SIZE),
				to_sfixed(-0.8346,1,L_SIZE),
				to_sfixed(-0.8345,1,L_SIZE),
				to_sfixed(-0.8343,1,L_SIZE),
				to_sfixed(-0.8342,1,L_SIZE),
				to_sfixed(-0.8341,1,L_SIZE),
				to_sfixed(-0.8340,1,L_SIZE),
				to_sfixed(-0.8339,1,L_SIZE),
				to_sfixed(-0.8338,1,L_SIZE),
				to_sfixed(-0.8337,1,L_SIZE),
				to_sfixed(-0.8336,1,L_SIZE),
				to_sfixed(-0.8335,1,L_SIZE),
				to_sfixed(-0.8333,1,L_SIZE),
				to_sfixed(-0.8332,1,L_SIZE),
				to_sfixed(-0.8331,1,L_SIZE),
				to_sfixed(-0.8330,1,L_SIZE),
				to_sfixed(-0.8329,1,L_SIZE),
				to_sfixed(-0.8328,1,L_SIZE),
				to_sfixed(-0.8327,1,L_SIZE),
				to_sfixed(-0.8326,1,L_SIZE),
				to_sfixed(-0.8324,1,L_SIZE),
				to_sfixed(-0.8323,1,L_SIZE),
				to_sfixed(-0.8322,1,L_SIZE),
				to_sfixed(-0.8321,1,L_SIZE),
				to_sfixed(-0.8320,1,L_SIZE),
				to_sfixed(-0.8319,1,L_SIZE),
				to_sfixed(-0.8318,1,L_SIZE),
				to_sfixed(-0.8317,1,L_SIZE),
				to_sfixed(-0.8315,1,L_SIZE),
				to_sfixed(-0.8314,1,L_SIZE),
				to_sfixed(-0.8313,1,L_SIZE),
				to_sfixed(-0.8312,1,L_SIZE),
				to_sfixed(-0.8311,1,L_SIZE),
				to_sfixed(-0.8310,1,L_SIZE),
				to_sfixed(-0.8309,1,L_SIZE),
				to_sfixed(-0.8307,1,L_SIZE),
				to_sfixed(-0.8306,1,L_SIZE),
				to_sfixed(-0.8305,1,L_SIZE),
				to_sfixed(-0.8304,1,L_SIZE),
				to_sfixed(-0.8303,1,L_SIZE),
				to_sfixed(-0.8302,1,L_SIZE),
				to_sfixed(-0.8301,1,L_SIZE),
				to_sfixed(-0.8300,1,L_SIZE),
				to_sfixed(-0.8298,1,L_SIZE),
				to_sfixed(-0.8297,1,L_SIZE),
				to_sfixed(-0.8296,1,L_SIZE),
				to_sfixed(-0.8295,1,L_SIZE),
				to_sfixed(-0.8294,1,L_SIZE),
				to_sfixed(-0.8293,1,L_SIZE),
				to_sfixed(-0.8292,1,L_SIZE),
				to_sfixed(-0.8290,1,L_SIZE),
				to_sfixed(-0.8289,1,L_SIZE),
				to_sfixed(-0.8288,1,L_SIZE),
				to_sfixed(-0.8287,1,L_SIZE),
				to_sfixed(-0.8286,1,L_SIZE),
				to_sfixed(-0.8285,1,L_SIZE),
				to_sfixed(-0.8284,1,L_SIZE),
				to_sfixed(-0.8282,1,L_SIZE),
				to_sfixed(-0.8281,1,L_SIZE),
				to_sfixed(-0.8280,1,L_SIZE),
				to_sfixed(-0.8279,1,L_SIZE),
				to_sfixed(-0.8278,1,L_SIZE),
				to_sfixed(-0.8277,1,L_SIZE),
				to_sfixed(-0.8275,1,L_SIZE),
				to_sfixed(-0.8274,1,L_SIZE),
				to_sfixed(-0.8273,1,L_SIZE),
				to_sfixed(-0.8272,1,L_SIZE),
				to_sfixed(-0.8271,1,L_SIZE),
				to_sfixed(-0.8270,1,L_SIZE),
				to_sfixed(-0.8269,1,L_SIZE),
				to_sfixed(-0.8267,1,L_SIZE),
				to_sfixed(-0.8266,1,L_SIZE),
				to_sfixed(-0.8265,1,L_SIZE),
				to_sfixed(-0.8264,1,L_SIZE),
				to_sfixed(-0.8263,1,L_SIZE),
				to_sfixed(-0.8262,1,L_SIZE),
				to_sfixed(-0.8260,1,L_SIZE),
				to_sfixed(-0.8259,1,L_SIZE),
				to_sfixed(-0.8258,1,L_SIZE),
				to_sfixed(-0.8257,1,L_SIZE),
				to_sfixed(-0.8256,1,L_SIZE),
				to_sfixed(-0.8255,1,L_SIZE),
				to_sfixed(-0.8253,1,L_SIZE),
				to_sfixed(-0.8252,1,L_SIZE),
				to_sfixed(-0.8251,1,L_SIZE),
				to_sfixed(-0.8250,1,L_SIZE),
				to_sfixed(-0.8249,1,L_SIZE),
				to_sfixed(-0.8248,1,L_SIZE),
				to_sfixed(-0.8246,1,L_SIZE),
				to_sfixed(-0.8245,1,L_SIZE),
				to_sfixed(-0.8244,1,L_SIZE),
				to_sfixed(-0.8243,1,L_SIZE),
				to_sfixed(-0.8242,1,L_SIZE),
				to_sfixed(-0.8241,1,L_SIZE),
				to_sfixed(-0.8239,1,L_SIZE),
				to_sfixed(-0.8238,1,L_SIZE),
				to_sfixed(-0.8237,1,L_SIZE),
				to_sfixed(-0.8236,1,L_SIZE),
				to_sfixed(-0.8235,1,L_SIZE),
				to_sfixed(-0.8233,1,L_SIZE),
				to_sfixed(-0.8232,1,L_SIZE),
				to_sfixed(-0.8231,1,L_SIZE),
				to_sfixed(-0.8230,1,L_SIZE),
				to_sfixed(-0.8229,1,L_SIZE),
				to_sfixed(-0.8228,1,L_SIZE),
				to_sfixed(-0.8226,1,L_SIZE),
				to_sfixed(-0.8225,1,L_SIZE),
				to_sfixed(-0.8224,1,L_SIZE),
				to_sfixed(-0.8223,1,L_SIZE),
				to_sfixed(-0.8222,1,L_SIZE),
				to_sfixed(-0.8220,1,L_SIZE),
				to_sfixed(-0.8219,1,L_SIZE),
				to_sfixed(-0.8218,1,L_SIZE),
				to_sfixed(-0.8217,1,L_SIZE),
				to_sfixed(-0.8216,1,L_SIZE),
				to_sfixed(-0.8214,1,L_SIZE),
				to_sfixed(-0.8213,1,L_SIZE),
				to_sfixed(-0.8212,1,L_SIZE),
				to_sfixed(-0.8211,1,L_SIZE),
				to_sfixed(-0.8210,1,L_SIZE),
				to_sfixed(-0.8209,1,L_SIZE),
				to_sfixed(-0.8207,1,L_SIZE),
				to_sfixed(-0.8206,1,L_SIZE),
				to_sfixed(-0.8205,1,L_SIZE),
				to_sfixed(-0.8204,1,L_SIZE),
				to_sfixed(-0.8203,1,L_SIZE),
				to_sfixed(-0.8201,1,L_SIZE),
				to_sfixed(-0.8200,1,L_SIZE),
				to_sfixed(-0.8199,1,L_SIZE),
				to_sfixed(-0.8198,1,L_SIZE),
				to_sfixed(-0.8197,1,L_SIZE),
				to_sfixed(-0.8195,1,L_SIZE),
				to_sfixed(-0.8194,1,L_SIZE),
				to_sfixed(-0.8193,1,L_SIZE),
				to_sfixed(-0.8192,1,L_SIZE),
				to_sfixed(-0.8191,1,L_SIZE),
				to_sfixed(-0.8189,1,L_SIZE),
				to_sfixed(-0.8188,1,L_SIZE),
				to_sfixed(-0.8187,1,L_SIZE),
				to_sfixed(-0.8186,1,L_SIZE),
				to_sfixed(-0.8184,1,L_SIZE),
				to_sfixed(-0.8183,1,L_SIZE),
				to_sfixed(-0.8182,1,L_SIZE),
				to_sfixed(-0.8181,1,L_SIZE),
				to_sfixed(-0.8180,1,L_SIZE),
				to_sfixed(-0.8178,1,L_SIZE),
				to_sfixed(-0.8177,1,L_SIZE),
				to_sfixed(-0.8176,1,L_SIZE),
				to_sfixed(-0.8175,1,L_SIZE),
				to_sfixed(-0.8174,1,L_SIZE),
				to_sfixed(-0.8172,1,L_SIZE),
				to_sfixed(-0.8171,1,L_SIZE),
				to_sfixed(-0.8170,1,L_SIZE),
				to_sfixed(-0.8169,1,L_SIZE),
				to_sfixed(-0.8167,1,L_SIZE),
				to_sfixed(-0.8166,1,L_SIZE),
				to_sfixed(-0.8165,1,L_SIZE),
				to_sfixed(-0.8164,1,L_SIZE),
				to_sfixed(-0.8163,1,L_SIZE),
				to_sfixed(-0.8161,1,L_SIZE),
				to_sfixed(-0.8160,1,L_SIZE),
				to_sfixed(-0.8159,1,L_SIZE),
				to_sfixed(-0.8158,1,L_SIZE),
				to_sfixed(-0.8156,1,L_SIZE),
				to_sfixed(-0.8155,1,L_SIZE),
				to_sfixed(-0.8154,1,L_SIZE),
				to_sfixed(-0.8153,1,L_SIZE),
				to_sfixed(-0.8152,1,L_SIZE),
				to_sfixed(-0.8150,1,L_SIZE),
				to_sfixed(-0.8149,1,L_SIZE),
				to_sfixed(-0.8148,1,L_SIZE),
				to_sfixed(-0.8147,1,L_SIZE),
				to_sfixed(-0.8145,1,L_SIZE),
				to_sfixed(-0.8144,1,L_SIZE),
				to_sfixed(-0.8143,1,L_SIZE),
				to_sfixed(-0.8142,1,L_SIZE),
				to_sfixed(-0.8140,1,L_SIZE),
				to_sfixed(-0.8139,1,L_SIZE),
				to_sfixed(-0.8138,1,L_SIZE),
				to_sfixed(-0.8137,1,L_SIZE),
				to_sfixed(-0.8136,1,L_SIZE),
				to_sfixed(-0.8134,1,L_SIZE),
				to_sfixed(-0.8133,1,L_SIZE),
				to_sfixed(-0.8132,1,L_SIZE),
				to_sfixed(-0.8131,1,L_SIZE),
				to_sfixed(-0.8129,1,L_SIZE),
				to_sfixed(-0.8128,1,L_SIZE),
				to_sfixed(-0.8127,1,L_SIZE),
				to_sfixed(-0.8126,1,L_SIZE),
				to_sfixed(-0.8124,1,L_SIZE),
				to_sfixed(-0.8123,1,L_SIZE),
				to_sfixed(-0.8122,1,L_SIZE),
				to_sfixed(-0.8121,1,L_SIZE),
				to_sfixed(-0.8119,1,L_SIZE),
				to_sfixed(-0.8118,1,L_SIZE),
				to_sfixed(-0.8117,1,L_SIZE),
				to_sfixed(-0.8116,1,L_SIZE),
				to_sfixed(-0.8114,1,L_SIZE),
				to_sfixed(-0.8113,1,L_SIZE),
				to_sfixed(-0.8112,1,L_SIZE),
				to_sfixed(-0.8111,1,L_SIZE),
				to_sfixed(-0.8109,1,L_SIZE),
				to_sfixed(-0.8108,1,L_SIZE),
				to_sfixed(-0.8107,1,L_SIZE),
				to_sfixed(-0.8106,1,L_SIZE),
				to_sfixed(-0.8104,1,L_SIZE),
				to_sfixed(-0.8103,1,L_SIZE),
				to_sfixed(-0.8102,1,L_SIZE),
				to_sfixed(-0.8101,1,L_SIZE),
				to_sfixed(-0.8099,1,L_SIZE),
				to_sfixed(-0.8098,1,L_SIZE),
				to_sfixed(-0.8097,1,L_SIZE),
				to_sfixed(-0.8096,1,L_SIZE),
				to_sfixed(-0.8094,1,L_SIZE),
				to_sfixed(-0.8093,1,L_SIZE),
				to_sfixed(-0.8092,1,L_SIZE),
				to_sfixed(-0.8090,1,L_SIZE),
				to_sfixed(-0.8089,1,L_SIZE),
				to_sfixed(-0.8088,1,L_SIZE),
				to_sfixed(-0.8087,1,L_SIZE),
				to_sfixed(-0.8085,1,L_SIZE),
				to_sfixed(-0.8084,1,L_SIZE),
				to_sfixed(-0.8083,1,L_SIZE),
				to_sfixed(-0.8082,1,L_SIZE),
				to_sfixed(-0.8080,1,L_SIZE),
				to_sfixed(-0.8079,1,L_SIZE),
				to_sfixed(-0.8078,1,L_SIZE),
				to_sfixed(-0.8077,1,L_SIZE),
				to_sfixed(-0.8075,1,L_SIZE),
				to_sfixed(-0.8074,1,L_SIZE),
				to_sfixed(-0.8073,1,L_SIZE),
				to_sfixed(-0.8071,1,L_SIZE),
				to_sfixed(-0.8070,1,L_SIZE),
				to_sfixed(-0.8069,1,L_SIZE),
				to_sfixed(-0.8068,1,L_SIZE),
				to_sfixed(-0.8066,1,L_SIZE),
				to_sfixed(-0.8065,1,L_SIZE),
				to_sfixed(-0.8064,1,L_SIZE),
				to_sfixed(-0.8062,1,L_SIZE),
				to_sfixed(-0.8061,1,L_SIZE),
				to_sfixed(-0.8060,1,L_SIZE),
				to_sfixed(-0.8059,1,L_SIZE),
				to_sfixed(-0.8057,1,L_SIZE),
				to_sfixed(-0.8056,1,L_SIZE),
				to_sfixed(-0.8055,1,L_SIZE),
				to_sfixed(-0.8053,1,L_SIZE),
				to_sfixed(-0.8052,1,L_SIZE),
				to_sfixed(-0.8051,1,L_SIZE),
				to_sfixed(-0.8050,1,L_SIZE),
				to_sfixed(-0.8048,1,L_SIZE),
				to_sfixed(-0.8047,1,L_SIZE),
				to_sfixed(-0.8046,1,L_SIZE),
				to_sfixed(-0.8044,1,L_SIZE),
				to_sfixed(-0.8043,1,L_SIZE),
				to_sfixed(-0.8042,1,L_SIZE),
				to_sfixed(-0.8041,1,L_SIZE),
				to_sfixed(-0.8039,1,L_SIZE),
				to_sfixed(-0.8038,1,L_SIZE),
				to_sfixed(-0.8037,1,L_SIZE),
				to_sfixed(-0.8035,1,L_SIZE),
				to_sfixed(-0.8034,1,L_SIZE),
				to_sfixed(-0.8033,1,L_SIZE),
				to_sfixed(-0.8031,1,L_SIZE),
				to_sfixed(-0.8030,1,L_SIZE),
				to_sfixed(-0.8029,1,L_SIZE),
				to_sfixed(-0.8028,1,L_SIZE),
				to_sfixed(-0.8026,1,L_SIZE),
				to_sfixed(-0.8025,1,L_SIZE),
				to_sfixed(-0.8024,1,L_SIZE),
				to_sfixed(-0.8022,1,L_SIZE),
				to_sfixed(-0.8021,1,L_SIZE),
				to_sfixed(-0.8020,1,L_SIZE),
				to_sfixed(-0.8018,1,L_SIZE),
				to_sfixed(-0.8017,1,L_SIZE),
				to_sfixed(-0.8016,1,L_SIZE),
				to_sfixed(-0.8015,1,L_SIZE),
				to_sfixed(-0.8013,1,L_SIZE),
				to_sfixed(-0.8012,1,L_SIZE),
				to_sfixed(-0.8011,1,L_SIZE),
				to_sfixed(-0.8009,1,L_SIZE),
				to_sfixed(-0.8008,1,L_SIZE),
				to_sfixed(-0.8007,1,L_SIZE),
				to_sfixed(-0.8005,1,L_SIZE),
				to_sfixed(-0.8004,1,L_SIZE),
				to_sfixed(-0.8003,1,L_SIZE),
				to_sfixed(-0.8001,1,L_SIZE),
				to_sfixed(-0.8000,1,L_SIZE),
				to_sfixed(-0.7999,1,L_SIZE),
				to_sfixed(-0.7997,1,L_SIZE),
				to_sfixed(-0.7996,1,L_SIZE),
				to_sfixed(-0.7995,1,L_SIZE),
				to_sfixed(-0.7993,1,L_SIZE),
				to_sfixed(-0.7992,1,L_SIZE),
				to_sfixed(-0.7991,1,L_SIZE),
				to_sfixed(-0.7990,1,L_SIZE),
				to_sfixed(-0.7988,1,L_SIZE),
				to_sfixed(-0.7987,1,L_SIZE),
				to_sfixed(-0.7986,1,L_SIZE),
				to_sfixed(-0.7984,1,L_SIZE),
				to_sfixed(-0.7983,1,L_SIZE),
				to_sfixed(-0.7982,1,L_SIZE),
				to_sfixed(-0.7980,1,L_SIZE),
				to_sfixed(-0.7979,1,L_SIZE),
				to_sfixed(-0.7978,1,L_SIZE),
				to_sfixed(-0.7976,1,L_SIZE),
				to_sfixed(-0.7975,1,L_SIZE),
				to_sfixed(-0.7974,1,L_SIZE),
				to_sfixed(-0.7972,1,L_SIZE),
				to_sfixed(-0.7971,1,L_SIZE),
				to_sfixed(-0.7970,1,L_SIZE),
				to_sfixed(-0.7968,1,L_SIZE),
				to_sfixed(-0.7967,1,L_SIZE),
				to_sfixed(-0.7966,1,L_SIZE),
				to_sfixed(-0.7964,1,L_SIZE),
				to_sfixed(-0.7963,1,L_SIZE),
				to_sfixed(-0.7962,1,L_SIZE),
				to_sfixed(-0.7960,1,L_SIZE),
				to_sfixed(-0.7959,1,L_SIZE),
				to_sfixed(-0.7957,1,L_SIZE),
				to_sfixed(-0.7956,1,L_SIZE),
				to_sfixed(-0.7955,1,L_SIZE),
				to_sfixed(-0.7953,1,L_SIZE),
				to_sfixed(-0.7952,1,L_SIZE),
				to_sfixed(-0.7951,1,L_SIZE),
				to_sfixed(-0.7949,1,L_SIZE),
				to_sfixed(-0.7948,1,L_SIZE),
				to_sfixed(-0.7947,1,L_SIZE),
				to_sfixed(-0.7945,1,L_SIZE),
				to_sfixed(-0.7944,1,L_SIZE),
				to_sfixed(-0.7943,1,L_SIZE),
				to_sfixed(-0.7941,1,L_SIZE),
				to_sfixed(-0.7940,1,L_SIZE),
				to_sfixed(-0.7939,1,L_SIZE),
				to_sfixed(-0.7937,1,L_SIZE),
				to_sfixed(-0.7936,1,L_SIZE),
				to_sfixed(-0.7935,1,L_SIZE),
				to_sfixed(-0.7933,1,L_SIZE),
				to_sfixed(-0.7932,1,L_SIZE),
				to_sfixed(-0.7930,1,L_SIZE),
				to_sfixed(-0.7929,1,L_SIZE),
				to_sfixed(-0.7928,1,L_SIZE),
				to_sfixed(-0.7926,1,L_SIZE),
				to_sfixed(-0.7925,1,L_SIZE),
				to_sfixed(-0.7924,1,L_SIZE),
				to_sfixed(-0.7922,1,L_SIZE),
				to_sfixed(-0.7921,1,L_SIZE),
				to_sfixed(-0.7920,1,L_SIZE),
				to_sfixed(-0.7918,1,L_SIZE),
				to_sfixed(-0.7917,1,L_SIZE),
				to_sfixed(-0.7915,1,L_SIZE),
				to_sfixed(-0.7914,1,L_SIZE),
				to_sfixed(-0.7913,1,L_SIZE),
				to_sfixed(-0.7911,1,L_SIZE),
				to_sfixed(-0.7910,1,L_SIZE),
				to_sfixed(-0.7909,1,L_SIZE),
				to_sfixed(-0.7907,1,L_SIZE),
				to_sfixed(-0.7906,1,L_SIZE),
				to_sfixed(-0.7905,1,L_SIZE),
				to_sfixed(-0.7903,1,L_SIZE),
				to_sfixed(-0.7902,1,L_SIZE),
				to_sfixed(-0.7900,1,L_SIZE),
				to_sfixed(-0.7899,1,L_SIZE),
				to_sfixed(-0.7898,1,L_SIZE),
				to_sfixed(-0.7896,1,L_SIZE),
				to_sfixed(-0.7895,1,L_SIZE),
				to_sfixed(-0.7893,1,L_SIZE),
				to_sfixed(-0.7892,1,L_SIZE),
				to_sfixed(-0.7891,1,L_SIZE),
				to_sfixed(-0.7889,1,L_SIZE),
				to_sfixed(-0.7888,1,L_SIZE),
				to_sfixed(-0.7887,1,L_SIZE),
				to_sfixed(-0.7885,1,L_SIZE),
				to_sfixed(-0.7884,1,L_SIZE),
				to_sfixed(-0.7882,1,L_SIZE),
				to_sfixed(-0.7881,1,L_SIZE),
				to_sfixed(-0.7880,1,L_SIZE),
				to_sfixed(-0.7878,1,L_SIZE),
				to_sfixed(-0.7877,1,L_SIZE),
				to_sfixed(-0.7875,1,L_SIZE),
				to_sfixed(-0.7874,1,L_SIZE),
				to_sfixed(-0.7873,1,L_SIZE),
				to_sfixed(-0.7871,1,L_SIZE),
				to_sfixed(-0.7870,1,L_SIZE),
				to_sfixed(-0.7869,1,L_SIZE),
				to_sfixed(-0.7867,1,L_SIZE),
				to_sfixed(-0.7866,1,L_SIZE),
				to_sfixed(-0.7864,1,L_SIZE),
				to_sfixed(-0.7863,1,L_SIZE),
				to_sfixed(-0.7862,1,L_SIZE),
				to_sfixed(-0.7860,1,L_SIZE),
				to_sfixed(-0.7859,1,L_SIZE),
				to_sfixed(-0.7857,1,L_SIZE),
				to_sfixed(-0.7856,1,L_SIZE),
				to_sfixed(-0.7855,1,L_SIZE),
				to_sfixed(-0.7853,1,L_SIZE),
				to_sfixed(-0.7852,1,L_SIZE),
				to_sfixed(-0.7850,1,L_SIZE),
				to_sfixed(-0.7849,1,L_SIZE),
				to_sfixed(-0.7848,1,L_SIZE),
				to_sfixed(-0.7846,1,L_SIZE),
				to_sfixed(-0.7845,1,L_SIZE),
				to_sfixed(-0.7843,1,L_SIZE),
				to_sfixed(-0.7842,1,L_SIZE),
				to_sfixed(-0.7840,1,L_SIZE),
				to_sfixed(-0.7839,1,L_SIZE),
				to_sfixed(-0.7838,1,L_SIZE),
				to_sfixed(-0.7836,1,L_SIZE),
				to_sfixed(-0.7835,1,L_SIZE),
				to_sfixed(-0.7833,1,L_SIZE),
				to_sfixed(-0.7832,1,L_SIZE),
				to_sfixed(-0.7831,1,L_SIZE),
				to_sfixed(-0.7829,1,L_SIZE),
				to_sfixed(-0.7828,1,L_SIZE),
				to_sfixed(-0.7826,1,L_SIZE),
				to_sfixed(-0.7825,1,L_SIZE),
				to_sfixed(-0.7823,1,L_SIZE),
				to_sfixed(-0.7822,1,L_SIZE),
				to_sfixed(-0.7821,1,L_SIZE),
				to_sfixed(-0.7819,1,L_SIZE),
				to_sfixed(-0.7818,1,L_SIZE),
				to_sfixed(-0.7816,1,L_SIZE),
				to_sfixed(-0.7815,1,L_SIZE),
				to_sfixed(-0.7814,1,L_SIZE),
				to_sfixed(-0.7812,1,L_SIZE),
				to_sfixed(-0.7811,1,L_SIZE),
				to_sfixed(-0.7809,1,L_SIZE),
				to_sfixed(-0.7808,1,L_SIZE),
				to_sfixed(-0.7806,1,L_SIZE),
				to_sfixed(-0.7805,1,L_SIZE),
				to_sfixed(-0.7803,1,L_SIZE),
				to_sfixed(-0.7802,1,L_SIZE),
				to_sfixed(-0.7801,1,L_SIZE),
				to_sfixed(-0.7799,1,L_SIZE),
				to_sfixed(-0.7798,1,L_SIZE),
				to_sfixed(-0.7796,1,L_SIZE),
				to_sfixed(-0.7795,1,L_SIZE),
				to_sfixed(-0.7793,1,L_SIZE),
				to_sfixed(-0.7792,1,L_SIZE),
				to_sfixed(-0.7791,1,L_SIZE),
				to_sfixed(-0.7789,1,L_SIZE),
				to_sfixed(-0.7788,1,L_SIZE),
				to_sfixed(-0.7786,1,L_SIZE),
				to_sfixed(-0.7785,1,L_SIZE),
				to_sfixed(-0.7783,1,L_SIZE),
				to_sfixed(-0.7782,1,L_SIZE),
				to_sfixed(-0.7780,1,L_SIZE),
				to_sfixed(-0.7779,1,L_SIZE),
				to_sfixed(-0.7778,1,L_SIZE),
				to_sfixed(-0.7776,1,L_SIZE),
				to_sfixed(-0.7775,1,L_SIZE),
				to_sfixed(-0.7773,1,L_SIZE),
				to_sfixed(-0.7772,1,L_SIZE),
				to_sfixed(-0.7770,1,L_SIZE),
				to_sfixed(-0.7769,1,L_SIZE),
				to_sfixed(-0.7767,1,L_SIZE),
				to_sfixed(-0.7766,1,L_SIZE),
				to_sfixed(-0.7765,1,L_SIZE),
				to_sfixed(-0.7763,1,L_SIZE),
				to_sfixed(-0.7762,1,L_SIZE),
				to_sfixed(-0.7760,1,L_SIZE),
				to_sfixed(-0.7759,1,L_SIZE),
				to_sfixed(-0.7757,1,L_SIZE),
				to_sfixed(-0.7756,1,L_SIZE),
				to_sfixed(-0.7754,1,L_SIZE),
				to_sfixed(-0.7753,1,L_SIZE),
				to_sfixed(-0.7751,1,L_SIZE),
				to_sfixed(-0.7750,1,L_SIZE),
				to_sfixed(-0.7748,1,L_SIZE),
				to_sfixed(-0.7747,1,L_SIZE),
				to_sfixed(-0.7746,1,L_SIZE),
				to_sfixed(-0.7744,1,L_SIZE),
				to_sfixed(-0.7743,1,L_SIZE),
				to_sfixed(-0.7741,1,L_SIZE),
				to_sfixed(-0.7740,1,L_SIZE),
				to_sfixed(-0.7738,1,L_SIZE),
				to_sfixed(-0.7737,1,L_SIZE),
				to_sfixed(-0.7735,1,L_SIZE),
				to_sfixed(-0.7734,1,L_SIZE),
				to_sfixed(-0.7732,1,L_SIZE),
				to_sfixed(-0.7731,1,L_SIZE),
				to_sfixed(-0.7729,1,L_SIZE),
				to_sfixed(-0.7728,1,L_SIZE),
				to_sfixed(-0.7726,1,L_SIZE),
				to_sfixed(-0.7725,1,L_SIZE),
				to_sfixed(-0.7723,1,L_SIZE),
				to_sfixed(-0.7722,1,L_SIZE),
				to_sfixed(-0.7721,1,L_SIZE),
				to_sfixed(-0.7719,1,L_SIZE),
				to_sfixed(-0.7718,1,L_SIZE),
				to_sfixed(-0.7716,1,L_SIZE),
				to_sfixed(-0.7715,1,L_SIZE),
				to_sfixed(-0.7713,1,L_SIZE),
				to_sfixed(-0.7712,1,L_SIZE),
				to_sfixed(-0.7710,1,L_SIZE),
				to_sfixed(-0.7709,1,L_SIZE),
				to_sfixed(-0.7707,1,L_SIZE),
				to_sfixed(-0.7706,1,L_SIZE),
				to_sfixed(-0.7704,1,L_SIZE),
				to_sfixed(-0.7703,1,L_SIZE),
				to_sfixed(-0.7701,1,L_SIZE),
				to_sfixed(-0.7700,1,L_SIZE),
				to_sfixed(-0.7698,1,L_SIZE),
				to_sfixed(-0.7697,1,L_SIZE),
				to_sfixed(-0.7695,1,L_SIZE),
				to_sfixed(-0.7694,1,L_SIZE),
				to_sfixed(-0.7692,1,L_SIZE),
				to_sfixed(-0.7691,1,L_SIZE),
				to_sfixed(-0.7689,1,L_SIZE),
				to_sfixed(-0.7688,1,L_SIZE),
				to_sfixed(-0.7686,1,L_SIZE),
				to_sfixed(-0.7685,1,L_SIZE),
				to_sfixed(-0.7683,1,L_SIZE),
				to_sfixed(-0.7682,1,L_SIZE),
				to_sfixed(-0.7680,1,L_SIZE),
				to_sfixed(-0.7679,1,L_SIZE),
				to_sfixed(-0.7677,1,L_SIZE),
				to_sfixed(-0.7676,1,L_SIZE),
				to_sfixed(-0.7674,1,L_SIZE),
				to_sfixed(-0.7673,1,L_SIZE),
				to_sfixed(-0.7671,1,L_SIZE),
				to_sfixed(-0.7670,1,L_SIZE),
				to_sfixed(-0.7668,1,L_SIZE),
				to_sfixed(-0.7667,1,L_SIZE),
				to_sfixed(-0.7665,1,L_SIZE),
				to_sfixed(-0.7664,1,L_SIZE),
				to_sfixed(-0.7662,1,L_SIZE),
				to_sfixed(-0.7661,1,L_SIZE),
				to_sfixed(-0.7659,1,L_SIZE),
				to_sfixed(-0.7658,1,L_SIZE),
				to_sfixed(-0.7656,1,L_SIZE),
				to_sfixed(-0.7655,1,L_SIZE),
				to_sfixed(-0.7653,1,L_SIZE),
				to_sfixed(-0.7652,1,L_SIZE),
				to_sfixed(-0.7650,1,L_SIZE),
				to_sfixed(-0.7649,1,L_SIZE),
				to_sfixed(-0.7647,1,L_SIZE),
				to_sfixed(-0.7646,1,L_SIZE),
				to_sfixed(-0.7644,1,L_SIZE),
				to_sfixed(-0.7642,1,L_SIZE),
				to_sfixed(-0.7641,1,L_SIZE),
				to_sfixed(-0.7639,1,L_SIZE),
				to_sfixed(-0.7638,1,L_SIZE),
				to_sfixed(-0.7636,1,L_SIZE),
				to_sfixed(-0.7635,1,L_SIZE),
				to_sfixed(-0.7633,1,L_SIZE),
				to_sfixed(-0.7632,1,L_SIZE),
				to_sfixed(-0.7630,1,L_SIZE),
				to_sfixed(-0.7629,1,L_SIZE),
				to_sfixed(-0.7627,1,L_SIZE),
				to_sfixed(-0.7626,1,L_SIZE),
				to_sfixed(-0.7624,1,L_SIZE),
				to_sfixed(-0.7623,1,L_SIZE),
				to_sfixed(-0.7621,1,L_SIZE),
				to_sfixed(-0.7620,1,L_SIZE),
				to_sfixed(-0.7618,1,L_SIZE),
				to_sfixed(-0.7616,1,L_SIZE),
				to_sfixed(-0.7615,1,L_SIZE),
				to_sfixed(-0.7613,1,L_SIZE),
				to_sfixed(-0.7612,1,L_SIZE),
				to_sfixed(-0.7610,1,L_SIZE),
				to_sfixed(-0.7609,1,L_SIZE),
				to_sfixed(-0.7607,1,L_SIZE),
				to_sfixed(-0.7606,1,L_SIZE),
				to_sfixed(-0.7604,1,L_SIZE),
				to_sfixed(-0.7603,1,L_SIZE),
				to_sfixed(-0.7601,1,L_SIZE),
				to_sfixed(-0.7599,1,L_SIZE),
				to_sfixed(-0.7598,1,L_SIZE),
				to_sfixed(-0.7596,1,L_SIZE),
				to_sfixed(-0.7595,1,L_SIZE),
				to_sfixed(-0.7593,1,L_SIZE),
				to_sfixed(-0.7592,1,L_SIZE),
				to_sfixed(-0.7590,1,L_SIZE),
				to_sfixed(-0.7589,1,L_SIZE),
				to_sfixed(-0.7587,1,L_SIZE),
				to_sfixed(-0.7586,1,L_SIZE),
				to_sfixed(-0.7584,1,L_SIZE),
				to_sfixed(-0.7582,1,L_SIZE),
				to_sfixed(-0.7581,1,L_SIZE),
				to_sfixed(-0.7579,1,L_SIZE),
				to_sfixed(-0.7578,1,L_SIZE),
				to_sfixed(-0.7576,1,L_SIZE),
				to_sfixed(-0.7575,1,L_SIZE),
				to_sfixed(-0.7573,1,L_SIZE),
				to_sfixed(-0.7571,1,L_SIZE),
				to_sfixed(-0.7570,1,L_SIZE),
				to_sfixed(-0.7568,1,L_SIZE),
				to_sfixed(-0.7567,1,L_SIZE),
				to_sfixed(-0.7565,1,L_SIZE),
				to_sfixed(-0.7564,1,L_SIZE),
				to_sfixed(-0.7562,1,L_SIZE),
				to_sfixed(-0.7561,1,L_SIZE),
				to_sfixed(-0.7559,1,L_SIZE),
				to_sfixed(-0.7557,1,L_SIZE),
				to_sfixed(-0.7556,1,L_SIZE),
				to_sfixed(-0.7554,1,L_SIZE),
				to_sfixed(-0.7553,1,L_SIZE),
				to_sfixed(-0.7551,1,L_SIZE),
				to_sfixed(-0.7550,1,L_SIZE),
				to_sfixed(-0.7548,1,L_SIZE),
				to_sfixed(-0.7546,1,L_SIZE),
				to_sfixed(-0.7545,1,L_SIZE),
				to_sfixed(-0.7543,1,L_SIZE),
				to_sfixed(-0.7542,1,L_SIZE),
				to_sfixed(-0.7540,1,L_SIZE),
				to_sfixed(-0.7538,1,L_SIZE),
				to_sfixed(-0.7537,1,L_SIZE),
				to_sfixed(-0.7535,1,L_SIZE),
				to_sfixed(-0.7534,1,L_SIZE),
				to_sfixed(-0.7532,1,L_SIZE),
				to_sfixed(-0.7531,1,L_SIZE),
				to_sfixed(-0.7529,1,L_SIZE),
				to_sfixed(-0.7527,1,L_SIZE),
				to_sfixed(-0.7526,1,L_SIZE),
				to_sfixed(-0.7524,1,L_SIZE),
				to_sfixed(-0.7523,1,L_SIZE),
				to_sfixed(-0.7521,1,L_SIZE),
				to_sfixed(-0.7519,1,L_SIZE),
				to_sfixed(-0.7518,1,L_SIZE),
				to_sfixed(-0.7516,1,L_SIZE),
				to_sfixed(-0.7515,1,L_SIZE),
				to_sfixed(-0.7513,1,L_SIZE),
				to_sfixed(-0.7511,1,L_SIZE),
				to_sfixed(-0.7510,1,L_SIZE),
				to_sfixed(-0.7508,1,L_SIZE),
				to_sfixed(-0.7507,1,L_SIZE),
				to_sfixed(-0.7505,1,L_SIZE),
				to_sfixed(-0.7503,1,L_SIZE),
				to_sfixed(-0.7502,1,L_SIZE),
				to_sfixed(-0.7500,1,L_SIZE),
				to_sfixed(-0.7499,1,L_SIZE),
				to_sfixed(-0.7497,1,L_SIZE),
				to_sfixed(-0.7495,1,L_SIZE),
				to_sfixed(-0.7494,1,L_SIZE),
				to_sfixed(-0.7492,1,L_SIZE),
				to_sfixed(-0.7491,1,L_SIZE),
				to_sfixed(-0.7489,1,L_SIZE),
				to_sfixed(-0.7487,1,L_SIZE),
				to_sfixed(-0.7486,1,L_SIZE),
				to_sfixed(-0.7484,1,L_SIZE),
				to_sfixed(-0.7483,1,L_SIZE),
				to_sfixed(-0.7481,1,L_SIZE),
				to_sfixed(-0.7479,1,L_SIZE),
				to_sfixed(-0.7478,1,L_SIZE),
				to_sfixed(-0.7476,1,L_SIZE),
				to_sfixed(-0.7475,1,L_SIZE),
				to_sfixed(-0.7473,1,L_SIZE),
				to_sfixed(-0.7471,1,L_SIZE),
				to_sfixed(-0.7470,1,L_SIZE),
				to_sfixed(-0.7468,1,L_SIZE),
				to_sfixed(-0.7466,1,L_SIZE),
				to_sfixed(-0.7465,1,L_SIZE),
				to_sfixed(-0.7463,1,L_SIZE),
				to_sfixed(-0.7462,1,L_SIZE),
				to_sfixed(-0.7460,1,L_SIZE),
				to_sfixed(-0.7458,1,L_SIZE),
				to_sfixed(-0.7457,1,L_SIZE),
				to_sfixed(-0.7455,1,L_SIZE),
				to_sfixed(-0.7453,1,L_SIZE),
				to_sfixed(-0.7452,1,L_SIZE),
				to_sfixed(-0.7450,1,L_SIZE),
				to_sfixed(-0.7449,1,L_SIZE),
				to_sfixed(-0.7447,1,L_SIZE),
				to_sfixed(-0.7445,1,L_SIZE),
				to_sfixed(-0.7444,1,L_SIZE),
				to_sfixed(-0.7442,1,L_SIZE),
				to_sfixed(-0.7440,1,L_SIZE),
				to_sfixed(-0.7439,1,L_SIZE),
				to_sfixed(-0.7437,1,L_SIZE),
				to_sfixed(-0.7436,1,L_SIZE),
				to_sfixed(-0.7434,1,L_SIZE),
				to_sfixed(-0.7432,1,L_SIZE),
				to_sfixed(-0.7431,1,L_SIZE),
				to_sfixed(-0.7429,1,L_SIZE),
				to_sfixed(-0.7427,1,L_SIZE),
				to_sfixed(-0.7426,1,L_SIZE),
				to_sfixed(-0.7424,1,L_SIZE),
				to_sfixed(-0.7422,1,L_SIZE),
				to_sfixed(-0.7421,1,L_SIZE),
				to_sfixed(-0.7419,1,L_SIZE),
				to_sfixed(-0.7417,1,L_SIZE),
				to_sfixed(-0.7416,1,L_SIZE),
				to_sfixed(-0.7414,1,L_SIZE),
				to_sfixed(-0.7412,1,L_SIZE),
				to_sfixed(-0.7411,1,L_SIZE),
				to_sfixed(-0.7409,1,L_SIZE),
				to_sfixed(-0.7408,1,L_SIZE),
				to_sfixed(-0.7406,1,L_SIZE),
				to_sfixed(-0.7404,1,L_SIZE),
				to_sfixed(-0.7403,1,L_SIZE),
				to_sfixed(-0.7401,1,L_SIZE),
				to_sfixed(-0.7399,1,L_SIZE),
				to_sfixed(-0.7398,1,L_SIZE),
				to_sfixed(-0.7396,1,L_SIZE),
				to_sfixed(-0.7394,1,L_SIZE),
				to_sfixed(-0.7393,1,L_SIZE),
				to_sfixed(-0.7391,1,L_SIZE),
				to_sfixed(-0.7389,1,L_SIZE),
				to_sfixed(-0.7388,1,L_SIZE),
				to_sfixed(-0.7386,1,L_SIZE),
				to_sfixed(-0.7384,1,L_SIZE),
				to_sfixed(-0.7383,1,L_SIZE),
				to_sfixed(-0.7381,1,L_SIZE),
				to_sfixed(-0.7379,1,L_SIZE),
				to_sfixed(-0.7378,1,L_SIZE),
				to_sfixed(-0.7376,1,L_SIZE),
				to_sfixed(-0.7374,1,L_SIZE),
				to_sfixed(-0.7373,1,L_SIZE),
				to_sfixed(-0.7371,1,L_SIZE),
				to_sfixed(-0.7369,1,L_SIZE),
				to_sfixed(-0.7368,1,L_SIZE),
				to_sfixed(-0.7366,1,L_SIZE),
				to_sfixed(-0.7364,1,L_SIZE),
				to_sfixed(-0.7363,1,L_SIZE),
				to_sfixed(-0.7361,1,L_SIZE),
				to_sfixed(-0.7359,1,L_SIZE),
				to_sfixed(-0.7358,1,L_SIZE),
				to_sfixed(-0.7356,1,L_SIZE),
				to_sfixed(-0.7354,1,L_SIZE),
				to_sfixed(-0.7353,1,L_SIZE),
				to_sfixed(-0.7351,1,L_SIZE),
				to_sfixed(-0.7349,1,L_SIZE),
				to_sfixed(-0.7347,1,L_SIZE),
				to_sfixed(-0.7346,1,L_SIZE),
				to_sfixed(-0.7344,1,L_SIZE),
				to_sfixed(-0.7342,1,L_SIZE),
				to_sfixed(-0.7341,1,L_SIZE),
				to_sfixed(-0.7339,1,L_SIZE),
				to_sfixed(-0.7337,1,L_SIZE),
				to_sfixed(-0.7336,1,L_SIZE),
				to_sfixed(-0.7334,1,L_SIZE),
				to_sfixed(-0.7332,1,L_SIZE),
				to_sfixed(-0.7331,1,L_SIZE),
				to_sfixed(-0.7329,1,L_SIZE),
				to_sfixed(-0.7327,1,L_SIZE),
				to_sfixed(-0.7325,1,L_SIZE),
				to_sfixed(-0.7324,1,L_SIZE),
				to_sfixed(-0.7322,1,L_SIZE),
				to_sfixed(-0.7320,1,L_SIZE),
				to_sfixed(-0.7319,1,L_SIZE),
				to_sfixed(-0.7317,1,L_SIZE),
				to_sfixed(-0.7315,1,L_SIZE),
				to_sfixed(-0.7314,1,L_SIZE),
				to_sfixed(-0.7312,1,L_SIZE),
				to_sfixed(-0.7310,1,L_SIZE),
				to_sfixed(-0.7308,1,L_SIZE),
				to_sfixed(-0.7307,1,L_SIZE),
				to_sfixed(-0.7305,1,L_SIZE),
				to_sfixed(-0.7303,1,L_SIZE),
				to_sfixed(-0.7302,1,L_SIZE),
				to_sfixed(-0.7300,1,L_SIZE),
				to_sfixed(-0.7298,1,L_SIZE),
				to_sfixed(-0.7297,1,L_SIZE),
				to_sfixed(-0.7295,1,L_SIZE),
				to_sfixed(-0.7293,1,L_SIZE),
				to_sfixed(-0.7291,1,L_SIZE),
				to_sfixed(-0.7290,1,L_SIZE),
				to_sfixed(-0.7288,1,L_SIZE),
				to_sfixed(-0.7286,1,L_SIZE),
				to_sfixed(-0.7284,1,L_SIZE),
				to_sfixed(-0.7283,1,L_SIZE),
				to_sfixed(-0.7281,1,L_SIZE),
				to_sfixed(-0.7279,1,L_SIZE),
				to_sfixed(-0.7278,1,L_SIZE),
				to_sfixed(-0.7276,1,L_SIZE),
				to_sfixed(-0.7274,1,L_SIZE),
				to_sfixed(-0.7272,1,L_SIZE),
				to_sfixed(-0.7271,1,L_SIZE),
				to_sfixed(-0.7269,1,L_SIZE),
				to_sfixed(-0.7267,1,L_SIZE),
				to_sfixed(-0.7266,1,L_SIZE),
				to_sfixed(-0.7264,1,L_SIZE),
				to_sfixed(-0.7262,1,L_SIZE),
				to_sfixed(-0.7260,1,L_SIZE),
				to_sfixed(-0.7259,1,L_SIZE),
				to_sfixed(-0.7257,1,L_SIZE),
				to_sfixed(-0.7255,1,L_SIZE),
				to_sfixed(-0.7253,1,L_SIZE),
				to_sfixed(-0.7252,1,L_SIZE),
				to_sfixed(-0.7250,1,L_SIZE),
				to_sfixed(-0.7248,1,L_SIZE),
				to_sfixed(-0.7246,1,L_SIZE),
				to_sfixed(-0.7245,1,L_SIZE),
				to_sfixed(-0.7243,1,L_SIZE),
				to_sfixed(-0.7241,1,L_SIZE),
				to_sfixed(-0.7239,1,L_SIZE),
				to_sfixed(-0.7238,1,L_SIZE),
				to_sfixed(-0.7236,1,L_SIZE),
				to_sfixed(-0.7234,1,L_SIZE),
				to_sfixed(-0.7233,1,L_SIZE),
				to_sfixed(-0.7231,1,L_SIZE),
				to_sfixed(-0.7229,1,L_SIZE),
				to_sfixed(-0.7227,1,L_SIZE),
				to_sfixed(-0.7226,1,L_SIZE),
				to_sfixed(-0.7224,1,L_SIZE),
				to_sfixed(-0.7222,1,L_SIZE),
				to_sfixed(-0.7220,1,L_SIZE),
				to_sfixed(-0.7219,1,L_SIZE),
				to_sfixed(-0.7217,1,L_SIZE),
				to_sfixed(-0.7215,1,L_SIZE),
				to_sfixed(-0.7213,1,L_SIZE),
				to_sfixed(-0.7211,1,L_SIZE),
				to_sfixed(-0.7210,1,L_SIZE),
				to_sfixed(-0.7208,1,L_SIZE),
				to_sfixed(-0.7206,1,L_SIZE),
				to_sfixed(-0.7204,1,L_SIZE),
				to_sfixed(-0.7203,1,L_SIZE),
				to_sfixed(-0.7201,1,L_SIZE),
				to_sfixed(-0.7199,1,L_SIZE),
				to_sfixed(-0.7197,1,L_SIZE),
				to_sfixed(-0.7196,1,L_SIZE),
				to_sfixed(-0.7194,1,L_SIZE),
				to_sfixed(-0.7192,1,L_SIZE),
				to_sfixed(-0.7190,1,L_SIZE),
				to_sfixed(-0.7189,1,L_SIZE),
				to_sfixed(-0.7187,1,L_SIZE),
				to_sfixed(-0.7185,1,L_SIZE),
				to_sfixed(-0.7183,1,L_SIZE),
				to_sfixed(-0.7181,1,L_SIZE),
				to_sfixed(-0.7180,1,L_SIZE),
				to_sfixed(-0.7178,1,L_SIZE),
				to_sfixed(-0.7176,1,L_SIZE),
				to_sfixed(-0.7174,1,L_SIZE),
				to_sfixed(-0.7173,1,L_SIZE),
				to_sfixed(-0.7171,1,L_SIZE),
				to_sfixed(-0.7169,1,L_SIZE),
				to_sfixed(-0.7167,1,L_SIZE),
				to_sfixed(-0.7165,1,L_SIZE),
				to_sfixed(-0.7164,1,L_SIZE),
				to_sfixed(-0.7162,1,L_SIZE),
				to_sfixed(-0.7160,1,L_SIZE),
				to_sfixed(-0.7158,1,L_SIZE),
				to_sfixed(-0.7157,1,L_SIZE),
				to_sfixed(-0.7155,1,L_SIZE),
				to_sfixed(-0.7153,1,L_SIZE),
				to_sfixed(-0.7151,1,L_SIZE),
				to_sfixed(-0.7149,1,L_SIZE),
				to_sfixed(-0.7148,1,L_SIZE),
				to_sfixed(-0.7146,1,L_SIZE),
				to_sfixed(-0.7144,1,L_SIZE),
				to_sfixed(-0.7142,1,L_SIZE),
				to_sfixed(-0.7140,1,L_SIZE),
				to_sfixed(-0.7139,1,L_SIZE),
				to_sfixed(-0.7137,1,L_SIZE),
				to_sfixed(-0.7135,1,L_SIZE),
				to_sfixed(-0.7133,1,L_SIZE),
				to_sfixed(-0.7131,1,L_SIZE),
				to_sfixed(-0.7130,1,L_SIZE),
				to_sfixed(-0.7128,1,L_SIZE),
				to_sfixed(-0.7126,1,L_SIZE),
				to_sfixed(-0.7124,1,L_SIZE),
				to_sfixed(-0.7122,1,L_SIZE),
				to_sfixed(-0.7121,1,L_SIZE),
				to_sfixed(-0.7119,1,L_SIZE),
				to_sfixed(-0.7117,1,L_SIZE),
				to_sfixed(-0.7115,1,L_SIZE),
				to_sfixed(-0.7113,1,L_SIZE),
				to_sfixed(-0.7112,1,L_SIZE),
				to_sfixed(-0.7110,1,L_SIZE),
				to_sfixed(-0.7108,1,L_SIZE),
				to_sfixed(-0.7106,1,L_SIZE),
				to_sfixed(-0.7104,1,L_SIZE),
				to_sfixed(-0.7103,1,L_SIZE),
				to_sfixed(-0.7101,1,L_SIZE),
				to_sfixed(-0.7099,1,L_SIZE),
				to_sfixed(-0.7097,1,L_SIZE),
				to_sfixed(-0.7095,1,L_SIZE),
				to_sfixed(-0.7093,1,L_SIZE),
				to_sfixed(-0.7092,1,L_SIZE),
				to_sfixed(-0.7090,1,L_SIZE),
				to_sfixed(-0.7088,1,L_SIZE),
				to_sfixed(-0.7086,1,L_SIZE),
				to_sfixed(-0.7084,1,L_SIZE),
				to_sfixed(-0.7083,1,L_SIZE),
				to_sfixed(-0.7081,1,L_SIZE),
				to_sfixed(-0.7079,1,L_SIZE),
				to_sfixed(-0.7077,1,L_SIZE),
				to_sfixed(-0.7075,1,L_SIZE),
				to_sfixed(-0.7073,1,L_SIZE),
				to_sfixed(-0.7072,1,L_SIZE),
				to_sfixed(-0.7070,1,L_SIZE),
				to_sfixed(-0.7068,1,L_SIZE),
				to_sfixed(-0.7066,1,L_SIZE),
				to_sfixed(-0.7064,1,L_SIZE),
				to_sfixed(-0.7062,1,L_SIZE),
				to_sfixed(-0.7061,1,L_SIZE),
				to_sfixed(-0.7059,1,L_SIZE),
				to_sfixed(-0.7057,1,L_SIZE),
				to_sfixed(-0.7055,1,L_SIZE),
				to_sfixed(-0.7053,1,L_SIZE),
				to_sfixed(-0.7051,1,L_SIZE),
				to_sfixed(-0.7050,1,L_SIZE),
				to_sfixed(-0.7048,1,L_SIZE),
				to_sfixed(-0.7046,1,L_SIZE),
				to_sfixed(-0.7044,1,L_SIZE),
				to_sfixed(-0.7042,1,L_SIZE),
				to_sfixed(-0.7040,1,L_SIZE),
				to_sfixed(-0.7038,1,L_SIZE),
				to_sfixed(-0.7037,1,L_SIZE),
				to_sfixed(-0.7035,1,L_SIZE),
				to_sfixed(-0.7033,1,L_SIZE),
				to_sfixed(-0.7031,1,L_SIZE),
				to_sfixed(-0.7029,1,L_SIZE),
				to_sfixed(-0.7027,1,L_SIZE),
				to_sfixed(-0.7025,1,L_SIZE),
				to_sfixed(-0.7024,1,L_SIZE),
				to_sfixed(-0.7022,1,L_SIZE),
				to_sfixed(-0.7020,1,L_SIZE),
				to_sfixed(-0.7018,1,L_SIZE),
				to_sfixed(-0.7016,1,L_SIZE),
				to_sfixed(-0.7014,1,L_SIZE),
				to_sfixed(-0.7012,1,L_SIZE),
				to_sfixed(-0.7011,1,L_SIZE),
				to_sfixed(-0.7009,1,L_SIZE),
				to_sfixed(-0.7007,1,L_SIZE),
				to_sfixed(-0.7005,1,L_SIZE),
				to_sfixed(-0.7003,1,L_SIZE),
				to_sfixed(-0.7001,1,L_SIZE),
				to_sfixed(-0.6999,1,L_SIZE),
				to_sfixed(-0.6998,1,L_SIZE),
				to_sfixed(-0.6996,1,L_SIZE),
				to_sfixed(-0.6994,1,L_SIZE),
				to_sfixed(-0.6992,1,L_SIZE),
				to_sfixed(-0.6990,1,L_SIZE),
				to_sfixed(-0.6988,1,L_SIZE),
				to_sfixed(-0.6986,1,L_SIZE),
				to_sfixed(-0.6984,1,L_SIZE),
				to_sfixed(-0.6983,1,L_SIZE),
				to_sfixed(-0.6981,1,L_SIZE),
				to_sfixed(-0.6979,1,L_SIZE),
				to_sfixed(-0.6977,1,L_SIZE),
				to_sfixed(-0.6975,1,L_SIZE),
				to_sfixed(-0.6973,1,L_SIZE),
				to_sfixed(-0.6971,1,L_SIZE),
				to_sfixed(-0.6969,1,L_SIZE),
				to_sfixed(-0.6968,1,L_SIZE),
				to_sfixed(-0.6966,1,L_SIZE),
				to_sfixed(-0.6964,1,L_SIZE),
				to_sfixed(-0.6962,1,L_SIZE),
				to_sfixed(-0.6960,1,L_SIZE),
				to_sfixed(-0.6958,1,L_SIZE),
				to_sfixed(-0.6956,1,L_SIZE),
				to_sfixed(-0.6954,1,L_SIZE),
				to_sfixed(-0.6952,1,L_SIZE),
				to_sfixed(-0.6951,1,L_SIZE),
				to_sfixed(-0.6949,1,L_SIZE),
				to_sfixed(-0.6947,1,L_SIZE),
				to_sfixed(-0.6945,1,L_SIZE),
				to_sfixed(-0.6943,1,L_SIZE),
				to_sfixed(-0.6941,1,L_SIZE),
				to_sfixed(-0.6939,1,L_SIZE),
				to_sfixed(-0.6937,1,L_SIZE),
				to_sfixed(-0.6935,1,L_SIZE),
				to_sfixed(-0.6933,1,L_SIZE),
				to_sfixed(-0.6932,1,L_SIZE),
				to_sfixed(-0.6930,1,L_SIZE),
				to_sfixed(-0.6928,1,L_SIZE),
				to_sfixed(-0.6926,1,L_SIZE),
				to_sfixed(-0.6924,1,L_SIZE),
				to_sfixed(-0.6922,1,L_SIZE),
				to_sfixed(-0.6920,1,L_SIZE),
				to_sfixed(-0.6918,1,L_SIZE),
				to_sfixed(-0.6916,1,L_SIZE),
				to_sfixed(-0.6914,1,L_SIZE),
				to_sfixed(-0.6912,1,L_SIZE),
				to_sfixed(-0.6911,1,L_SIZE),
				to_sfixed(-0.6909,1,L_SIZE),
				to_sfixed(-0.6907,1,L_SIZE),
				to_sfixed(-0.6905,1,L_SIZE),
				to_sfixed(-0.6903,1,L_SIZE),
				to_sfixed(-0.6901,1,L_SIZE),
				to_sfixed(-0.6899,1,L_SIZE),
				to_sfixed(-0.6897,1,L_SIZE),
				to_sfixed(-0.6895,1,L_SIZE),
				to_sfixed(-0.6893,1,L_SIZE),
				to_sfixed(-0.6891,1,L_SIZE),
				to_sfixed(-0.6889,1,L_SIZE),
				to_sfixed(-0.6888,1,L_SIZE),
				to_sfixed(-0.6886,1,L_SIZE),
				to_sfixed(-0.6884,1,L_SIZE),
				to_sfixed(-0.6882,1,L_SIZE),
				to_sfixed(-0.6880,1,L_SIZE),
				to_sfixed(-0.6878,1,L_SIZE),
				to_sfixed(-0.6876,1,L_SIZE),
				to_sfixed(-0.6874,1,L_SIZE),
				to_sfixed(-0.6872,1,L_SIZE),
				to_sfixed(-0.6870,1,L_SIZE),
				to_sfixed(-0.6868,1,L_SIZE),
				to_sfixed(-0.6866,1,L_SIZE),
				to_sfixed(-0.6864,1,L_SIZE),
				to_sfixed(-0.6862,1,L_SIZE),
				to_sfixed(-0.6860,1,L_SIZE),
				to_sfixed(-0.6859,1,L_SIZE),
				to_sfixed(-0.6857,1,L_SIZE),
				to_sfixed(-0.6855,1,L_SIZE),
				to_sfixed(-0.6853,1,L_SIZE),
				to_sfixed(-0.6851,1,L_SIZE),
				to_sfixed(-0.6849,1,L_SIZE),
				to_sfixed(-0.6847,1,L_SIZE),
				to_sfixed(-0.6845,1,L_SIZE),
				to_sfixed(-0.6843,1,L_SIZE),
				to_sfixed(-0.6841,1,L_SIZE),
				to_sfixed(-0.6839,1,L_SIZE),
				to_sfixed(-0.6837,1,L_SIZE),
				to_sfixed(-0.6835,1,L_SIZE),
				to_sfixed(-0.6833,1,L_SIZE),
				to_sfixed(-0.6831,1,L_SIZE),
				to_sfixed(-0.6829,1,L_SIZE),
				to_sfixed(-0.6827,1,L_SIZE),
				to_sfixed(-0.6825,1,L_SIZE),
				to_sfixed(-0.6823,1,L_SIZE),
				to_sfixed(-0.6822,1,L_SIZE),
				to_sfixed(-0.6820,1,L_SIZE),
				to_sfixed(-0.6818,1,L_SIZE),
				to_sfixed(-0.6816,1,L_SIZE),
				to_sfixed(-0.6814,1,L_SIZE),
				to_sfixed(-0.6812,1,L_SIZE),
				to_sfixed(-0.6810,1,L_SIZE),
				to_sfixed(-0.6808,1,L_SIZE),
				to_sfixed(-0.6806,1,L_SIZE),
				to_sfixed(-0.6804,1,L_SIZE),
				to_sfixed(-0.6802,1,L_SIZE),
				to_sfixed(-0.6800,1,L_SIZE),
				to_sfixed(-0.6798,1,L_SIZE),
				to_sfixed(-0.6796,1,L_SIZE),
				to_sfixed(-0.6794,1,L_SIZE),
				to_sfixed(-0.6792,1,L_SIZE),
				to_sfixed(-0.6790,1,L_SIZE),
				to_sfixed(-0.6788,1,L_SIZE),
				to_sfixed(-0.6786,1,L_SIZE),
				to_sfixed(-0.6784,1,L_SIZE),
				to_sfixed(-0.6782,1,L_SIZE),
				to_sfixed(-0.6780,1,L_SIZE),
				to_sfixed(-0.6778,1,L_SIZE),
				to_sfixed(-0.6776,1,L_SIZE),
				to_sfixed(-0.6774,1,L_SIZE),
				to_sfixed(-0.6772,1,L_SIZE),
				to_sfixed(-0.6770,1,L_SIZE),
				to_sfixed(-0.6768,1,L_SIZE),
				to_sfixed(-0.6766,1,L_SIZE),
				to_sfixed(-0.6764,1,L_SIZE),
				to_sfixed(-0.6762,1,L_SIZE),
				to_sfixed(-0.6760,1,L_SIZE),
				to_sfixed(-0.6758,1,L_SIZE),
				to_sfixed(-0.6756,1,L_SIZE),
				to_sfixed(-0.6754,1,L_SIZE),
				to_sfixed(-0.6752,1,L_SIZE),
				to_sfixed(-0.6750,1,L_SIZE),
				to_sfixed(-0.6748,1,L_SIZE),
				to_sfixed(-0.6746,1,L_SIZE),
				to_sfixed(-0.6744,1,L_SIZE),
				to_sfixed(-0.6742,1,L_SIZE),
				to_sfixed(-0.6740,1,L_SIZE),
				to_sfixed(-0.6738,1,L_SIZE),
				to_sfixed(-0.6736,1,L_SIZE),
				to_sfixed(-0.6734,1,L_SIZE),
				to_sfixed(-0.6732,1,L_SIZE),
				to_sfixed(-0.6730,1,L_SIZE),
				to_sfixed(-0.6728,1,L_SIZE),
				to_sfixed(-0.6726,1,L_SIZE),
				to_sfixed(-0.6724,1,L_SIZE),
				to_sfixed(-0.6722,1,L_SIZE),
				to_sfixed(-0.6720,1,L_SIZE),
				to_sfixed(-0.6718,1,L_SIZE),
				to_sfixed(-0.6716,1,L_SIZE),
				to_sfixed(-0.6714,1,L_SIZE),
				to_sfixed(-0.6712,1,L_SIZE),
				to_sfixed(-0.6710,1,L_SIZE),
				to_sfixed(-0.6708,1,L_SIZE),
				to_sfixed(-0.6706,1,L_SIZE),
				to_sfixed(-0.6704,1,L_SIZE),
				to_sfixed(-0.6702,1,L_SIZE),
				to_sfixed(-0.6700,1,L_SIZE),
				to_sfixed(-0.6698,1,L_SIZE),
				to_sfixed(-0.6696,1,L_SIZE),
				to_sfixed(-0.6694,1,L_SIZE),
				to_sfixed(-0.6692,1,L_SIZE),
				to_sfixed(-0.6690,1,L_SIZE),
				to_sfixed(-0.6688,1,L_SIZE),
				to_sfixed(-0.6686,1,L_SIZE),
				to_sfixed(-0.6684,1,L_SIZE),
				to_sfixed(-0.6682,1,L_SIZE),
				to_sfixed(-0.6680,1,L_SIZE),
				to_sfixed(-0.6678,1,L_SIZE),
				to_sfixed(-0.6676,1,L_SIZE),
				to_sfixed(-0.6674,1,L_SIZE),
				to_sfixed(-0.6672,1,L_SIZE),
				to_sfixed(-0.6670,1,L_SIZE),
				to_sfixed(-0.6668,1,L_SIZE),
				to_sfixed(-0.6666,1,L_SIZE),
				to_sfixed(-0.6664,1,L_SIZE),
				to_sfixed(-0.6662,1,L_SIZE),
				to_sfixed(-0.6660,1,L_SIZE),
				to_sfixed(-0.6658,1,L_SIZE),
				to_sfixed(-0.6656,1,L_SIZE),
				to_sfixed(-0.6654,1,L_SIZE),
				to_sfixed(-0.6652,1,L_SIZE),
				to_sfixed(-0.6650,1,L_SIZE),
				to_sfixed(-0.6647,1,L_SIZE),
				to_sfixed(-0.6645,1,L_SIZE),
				to_sfixed(-0.6643,1,L_SIZE),
				to_sfixed(-0.6641,1,L_SIZE),
				to_sfixed(-0.6639,1,L_SIZE),
				to_sfixed(-0.6637,1,L_SIZE),
				to_sfixed(-0.6635,1,L_SIZE),
				to_sfixed(-0.6633,1,L_SIZE),
				to_sfixed(-0.6631,1,L_SIZE),
				to_sfixed(-0.6629,1,L_SIZE),
				to_sfixed(-0.6627,1,L_SIZE),
				to_sfixed(-0.6625,1,L_SIZE),
				to_sfixed(-0.6623,1,L_SIZE),
				to_sfixed(-0.6621,1,L_SIZE),
				to_sfixed(-0.6619,1,L_SIZE),
				to_sfixed(-0.6617,1,L_SIZE),
				to_sfixed(-0.6615,1,L_SIZE),
				to_sfixed(-0.6613,1,L_SIZE),
				to_sfixed(-0.6611,1,L_SIZE),
				to_sfixed(-0.6608,1,L_SIZE),
				to_sfixed(-0.6606,1,L_SIZE),
				to_sfixed(-0.6604,1,L_SIZE),
				to_sfixed(-0.6602,1,L_SIZE),
				to_sfixed(-0.6600,1,L_SIZE),
				to_sfixed(-0.6598,1,L_SIZE),
				to_sfixed(-0.6596,1,L_SIZE),
				to_sfixed(-0.6594,1,L_SIZE),
				to_sfixed(-0.6592,1,L_SIZE),
				to_sfixed(-0.6590,1,L_SIZE),
				to_sfixed(-0.6588,1,L_SIZE),
				to_sfixed(-0.6586,1,L_SIZE),
				to_sfixed(-0.6584,1,L_SIZE),
				to_sfixed(-0.6582,1,L_SIZE),
				to_sfixed(-0.6579,1,L_SIZE),
				to_sfixed(-0.6577,1,L_SIZE),
				to_sfixed(-0.6575,1,L_SIZE),
				to_sfixed(-0.6573,1,L_SIZE),
				to_sfixed(-0.6571,1,L_SIZE),
				to_sfixed(-0.6569,1,L_SIZE),
				to_sfixed(-0.6567,1,L_SIZE),
				to_sfixed(-0.6565,1,L_SIZE),
				to_sfixed(-0.6563,1,L_SIZE),
				to_sfixed(-0.6561,1,L_SIZE),
				to_sfixed(-0.6559,1,L_SIZE),
				to_sfixed(-0.6557,1,L_SIZE),
				to_sfixed(-0.6554,1,L_SIZE),
				to_sfixed(-0.6552,1,L_SIZE),
				to_sfixed(-0.6550,1,L_SIZE),
				to_sfixed(-0.6548,1,L_SIZE),
				to_sfixed(-0.6546,1,L_SIZE),
				to_sfixed(-0.6544,1,L_SIZE),
				to_sfixed(-0.6542,1,L_SIZE),
				to_sfixed(-0.6540,1,L_SIZE),
				to_sfixed(-0.6538,1,L_SIZE),
				to_sfixed(-0.6536,1,L_SIZE),
				to_sfixed(-0.6534,1,L_SIZE),
				to_sfixed(-0.6531,1,L_SIZE),
				to_sfixed(-0.6529,1,L_SIZE),
				to_sfixed(-0.6527,1,L_SIZE),
				to_sfixed(-0.6525,1,L_SIZE),
				to_sfixed(-0.6523,1,L_SIZE),
				to_sfixed(-0.6521,1,L_SIZE),
				to_sfixed(-0.6519,1,L_SIZE),
				to_sfixed(-0.6517,1,L_SIZE),
				to_sfixed(-0.6515,1,L_SIZE),
				to_sfixed(-0.6512,1,L_SIZE),
				to_sfixed(-0.6510,1,L_SIZE),
				to_sfixed(-0.6508,1,L_SIZE),
				to_sfixed(-0.6506,1,L_SIZE),
				to_sfixed(-0.6504,1,L_SIZE),
				to_sfixed(-0.6502,1,L_SIZE),
				to_sfixed(-0.6500,1,L_SIZE),
				to_sfixed(-0.6498,1,L_SIZE),
				to_sfixed(-0.6496,1,L_SIZE),
				to_sfixed(-0.6493,1,L_SIZE),
				to_sfixed(-0.6491,1,L_SIZE),
				to_sfixed(-0.6489,1,L_SIZE),
				to_sfixed(-0.6487,1,L_SIZE),
				to_sfixed(-0.6485,1,L_SIZE),
				to_sfixed(-0.6483,1,L_SIZE),
				to_sfixed(-0.6481,1,L_SIZE),
				to_sfixed(-0.6479,1,L_SIZE),
				to_sfixed(-0.6477,1,L_SIZE),
				to_sfixed(-0.6474,1,L_SIZE),
				to_sfixed(-0.6472,1,L_SIZE),
				to_sfixed(-0.6470,1,L_SIZE),
				to_sfixed(-0.6468,1,L_SIZE),
				to_sfixed(-0.6466,1,L_SIZE),
				to_sfixed(-0.6464,1,L_SIZE),
				to_sfixed(-0.6462,1,L_SIZE),
				to_sfixed(-0.6459,1,L_SIZE),
				to_sfixed(-0.6457,1,L_SIZE),
				to_sfixed(-0.6455,1,L_SIZE),
				to_sfixed(-0.6453,1,L_SIZE),
				to_sfixed(-0.6451,1,L_SIZE),
				to_sfixed(-0.6449,1,L_SIZE),
				to_sfixed(-0.6447,1,L_SIZE),
				to_sfixed(-0.6444,1,L_SIZE),
				to_sfixed(-0.6442,1,L_SIZE),
				to_sfixed(-0.6440,1,L_SIZE),
				to_sfixed(-0.6438,1,L_SIZE),
				to_sfixed(-0.6436,1,L_SIZE),
				to_sfixed(-0.6434,1,L_SIZE),
				to_sfixed(-0.6432,1,L_SIZE),
				to_sfixed(-0.6429,1,L_SIZE),
				to_sfixed(-0.6427,1,L_SIZE),
				to_sfixed(-0.6425,1,L_SIZE),
				to_sfixed(-0.6423,1,L_SIZE),
				to_sfixed(-0.6421,1,L_SIZE),
				to_sfixed(-0.6419,1,L_SIZE),
				to_sfixed(-0.6417,1,L_SIZE),
				to_sfixed(-0.6414,1,L_SIZE),
				to_sfixed(-0.6412,1,L_SIZE),
				to_sfixed(-0.6410,1,L_SIZE),
				to_sfixed(-0.6408,1,L_SIZE),
				to_sfixed(-0.6406,1,L_SIZE),
				to_sfixed(-0.6404,1,L_SIZE),
				to_sfixed(-0.6401,1,L_SIZE),
				to_sfixed(-0.6399,1,L_SIZE),
				to_sfixed(-0.6397,1,L_SIZE),
				to_sfixed(-0.6395,1,L_SIZE),
				to_sfixed(-0.6393,1,L_SIZE),
				to_sfixed(-0.6391,1,L_SIZE),
				to_sfixed(-0.6388,1,L_SIZE),
				to_sfixed(-0.6386,1,L_SIZE),
				to_sfixed(-0.6384,1,L_SIZE),
				to_sfixed(-0.6382,1,L_SIZE),
				to_sfixed(-0.6380,1,L_SIZE),
				to_sfixed(-0.6378,1,L_SIZE),
				to_sfixed(-0.6375,1,L_SIZE),
				to_sfixed(-0.6373,1,L_SIZE),
				to_sfixed(-0.6371,1,L_SIZE),
				to_sfixed(-0.6369,1,L_SIZE),
				to_sfixed(-0.6367,1,L_SIZE),
				to_sfixed(-0.6365,1,L_SIZE),
				to_sfixed(-0.6362,1,L_SIZE),
				to_sfixed(-0.6360,1,L_SIZE),
				to_sfixed(-0.6358,1,L_SIZE),
				to_sfixed(-0.6356,1,L_SIZE),
				to_sfixed(-0.6354,1,L_SIZE),
				to_sfixed(-0.6351,1,L_SIZE),
				to_sfixed(-0.6349,1,L_SIZE),
				to_sfixed(-0.6347,1,L_SIZE),
				to_sfixed(-0.6345,1,L_SIZE),
				to_sfixed(-0.6343,1,L_SIZE),
				to_sfixed(-0.6341,1,L_SIZE),
				to_sfixed(-0.6338,1,L_SIZE),
				to_sfixed(-0.6336,1,L_SIZE),
				to_sfixed(-0.6334,1,L_SIZE),
				to_sfixed(-0.6332,1,L_SIZE),
				to_sfixed(-0.6330,1,L_SIZE),
				to_sfixed(-0.6327,1,L_SIZE),
				to_sfixed(-0.6325,1,L_SIZE),
				to_sfixed(-0.6323,1,L_SIZE),
				to_sfixed(-0.6321,1,L_SIZE),
				to_sfixed(-0.6319,1,L_SIZE),
				to_sfixed(-0.6316,1,L_SIZE),
				to_sfixed(-0.6314,1,L_SIZE),
				to_sfixed(-0.6312,1,L_SIZE),
				to_sfixed(-0.6310,1,L_SIZE),
				to_sfixed(-0.6308,1,L_SIZE),
				to_sfixed(-0.6305,1,L_SIZE),
				to_sfixed(-0.6303,1,L_SIZE),
				to_sfixed(-0.6301,1,L_SIZE),
				to_sfixed(-0.6299,1,L_SIZE),
				to_sfixed(-0.6297,1,L_SIZE),
				to_sfixed(-0.6294,1,L_SIZE),
				to_sfixed(-0.6292,1,L_SIZE),
				to_sfixed(-0.6290,1,L_SIZE),
				to_sfixed(-0.6288,1,L_SIZE),
				to_sfixed(-0.6285,1,L_SIZE),
				to_sfixed(-0.6283,1,L_SIZE),
				to_sfixed(-0.6281,1,L_SIZE),
				to_sfixed(-0.6279,1,L_SIZE),
				to_sfixed(-0.6277,1,L_SIZE),
				to_sfixed(-0.6274,1,L_SIZE),
				to_sfixed(-0.6272,1,L_SIZE),
				to_sfixed(-0.6270,1,L_SIZE),
				to_sfixed(-0.6268,1,L_SIZE),
				to_sfixed(-0.6266,1,L_SIZE),
				to_sfixed(-0.6263,1,L_SIZE),
				to_sfixed(-0.6261,1,L_SIZE),
				to_sfixed(-0.6259,1,L_SIZE),
				to_sfixed(-0.6257,1,L_SIZE),
				to_sfixed(-0.6254,1,L_SIZE),
				to_sfixed(-0.6252,1,L_SIZE),
				to_sfixed(-0.6250,1,L_SIZE),
				to_sfixed(-0.6248,1,L_SIZE),
				to_sfixed(-0.6245,1,L_SIZE),
				to_sfixed(-0.6243,1,L_SIZE),
				to_sfixed(-0.6241,1,L_SIZE),
				to_sfixed(-0.6239,1,L_SIZE),
				to_sfixed(-0.6237,1,L_SIZE),
				to_sfixed(-0.6234,1,L_SIZE),
				to_sfixed(-0.6232,1,L_SIZE),
				to_sfixed(-0.6230,1,L_SIZE),
				to_sfixed(-0.6228,1,L_SIZE),
				to_sfixed(-0.6225,1,L_SIZE),
				to_sfixed(-0.6223,1,L_SIZE),
				to_sfixed(-0.6221,1,L_SIZE),
				to_sfixed(-0.6219,1,L_SIZE),
				to_sfixed(-0.6216,1,L_SIZE),
				to_sfixed(-0.6214,1,L_SIZE),
				to_sfixed(-0.6212,1,L_SIZE),
				to_sfixed(-0.6210,1,L_SIZE),
				to_sfixed(-0.6207,1,L_SIZE),
				to_sfixed(-0.6205,1,L_SIZE),
				to_sfixed(-0.6203,1,L_SIZE),
				to_sfixed(-0.6201,1,L_SIZE),
				to_sfixed(-0.6198,1,L_SIZE),
				to_sfixed(-0.6196,1,L_SIZE),
				to_sfixed(-0.6194,1,L_SIZE),
				to_sfixed(-0.6192,1,L_SIZE),
				to_sfixed(-0.6189,1,L_SIZE),
				to_sfixed(-0.6187,1,L_SIZE),
				to_sfixed(-0.6185,1,L_SIZE),
				to_sfixed(-0.6183,1,L_SIZE),
				to_sfixed(-0.6180,1,L_SIZE),
				to_sfixed(-0.6178,1,L_SIZE),
				to_sfixed(-0.6176,1,L_SIZE),
				to_sfixed(-0.6173,1,L_SIZE),
				to_sfixed(-0.6171,1,L_SIZE),
				to_sfixed(-0.6169,1,L_SIZE),
				to_sfixed(-0.6167,1,L_SIZE),
				to_sfixed(-0.6164,1,L_SIZE),
				to_sfixed(-0.6162,1,L_SIZE),
				to_sfixed(-0.6160,1,L_SIZE),
				to_sfixed(-0.6158,1,L_SIZE),
				to_sfixed(-0.6155,1,L_SIZE),
				to_sfixed(-0.6153,1,L_SIZE),
				to_sfixed(-0.6151,1,L_SIZE),
				to_sfixed(-0.6148,1,L_SIZE),
				to_sfixed(-0.6146,1,L_SIZE),
				to_sfixed(-0.6144,1,L_SIZE),
				to_sfixed(-0.6142,1,L_SIZE),
				to_sfixed(-0.6139,1,L_SIZE),
				to_sfixed(-0.6137,1,L_SIZE),
				to_sfixed(-0.6135,1,L_SIZE),
				to_sfixed(-0.6132,1,L_SIZE),
				to_sfixed(-0.6130,1,L_SIZE),
				to_sfixed(-0.6128,1,L_SIZE),
				to_sfixed(-0.6126,1,L_SIZE),
				to_sfixed(-0.6123,1,L_SIZE),
				to_sfixed(-0.6121,1,L_SIZE),
				to_sfixed(-0.6119,1,L_SIZE),
				to_sfixed(-0.6116,1,L_SIZE),
				to_sfixed(-0.6114,1,L_SIZE),
				to_sfixed(-0.6112,1,L_SIZE),
				to_sfixed(-0.6110,1,L_SIZE),
				to_sfixed(-0.6107,1,L_SIZE),
				to_sfixed(-0.6105,1,L_SIZE),
				to_sfixed(-0.6103,1,L_SIZE),
				to_sfixed(-0.6100,1,L_SIZE),
				to_sfixed(-0.6098,1,L_SIZE),
				to_sfixed(-0.6096,1,L_SIZE),
				to_sfixed(-0.6093,1,L_SIZE),
				to_sfixed(-0.6091,1,L_SIZE),
				to_sfixed(-0.6089,1,L_SIZE),
				to_sfixed(-0.6087,1,L_SIZE),
				to_sfixed(-0.6084,1,L_SIZE),
				to_sfixed(-0.6082,1,L_SIZE),
				to_sfixed(-0.6080,1,L_SIZE),
				to_sfixed(-0.6077,1,L_SIZE),
				to_sfixed(-0.6075,1,L_SIZE),
				to_sfixed(-0.6073,1,L_SIZE),
				to_sfixed(-0.6070,1,L_SIZE),
				to_sfixed(-0.6068,1,L_SIZE),
				to_sfixed(-0.6066,1,L_SIZE),
				to_sfixed(-0.6063,1,L_SIZE),
				to_sfixed(-0.6061,1,L_SIZE),
				to_sfixed(-0.6059,1,L_SIZE),
				to_sfixed(-0.6057,1,L_SIZE),
				to_sfixed(-0.6054,1,L_SIZE),
				to_sfixed(-0.6052,1,L_SIZE),
				to_sfixed(-0.6050,1,L_SIZE),
				to_sfixed(-0.6047,1,L_SIZE),
				to_sfixed(-0.6045,1,L_SIZE),
				to_sfixed(-0.6043,1,L_SIZE),
				to_sfixed(-0.6040,1,L_SIZE),
				to_sfixed(-0.6038,1,L_SIZE),
				to_sfixed(-0.6036,1,L_SIZE),
				to_sfixed(-0.6033,1,L_SIZE),
				to_sfixed(-0.6031,1,L_SIZE),
				to_sfixed(-0.6029,1,L_SIZE),
				to_sfixed(-0.6026,1,L_SIZE),
				to_sfixed(-0.6024,1,L_SIZE),
				to_sfixed(-0.6022,1,L_SIZE),
				to_sfixed(-0.6019,1,L_SIZE),
				to_sfixed(-0.6017,1,L_SIZE),
				to_sfixed(-0.6015,1,L_SIZE),
				to_sfixed(-0.6012,1,L_SIZE),
				to_sfixed(-0.6010,1,L_SIZE),
				to_sfixed(-0.6008,1,L_SIZE),
				to_sfixed(-0.6005,1,L_SIZE),
				to_sfixed(-0.6003,1,L_SIZE),
				to_sfixed(-0.6001,1,L_SIZE),
				to_sfixed(-0.5998,1,L_SIZE),
				to_sfixed(-0.5996,1,L_SIZE),
				to_sfixed(-0.5994,1,L_SIZE),
				to_sfixed(-0.5991,1,L_SIZE),
				to_sfixed(-0.5989,1,L_SIZE),
				to_sfixed(-0.5986,1,L_SIZE),
				to_sfixed(-0.5984,1,L_SIZE),
				to_sfixed(-0.5982,1,L_SIZE),
				to_sfixed(-0.5979,1,L_SIZE),
				to_sfixed(-0.5977,1,L_SIZE),
				to_sfixed(-0.5975,1,L_SIZE),
				to_sfixed(-0.5972,1,L_SIZE),
				to_sfixed(-0.5970,1,L_SIZE),
				to_sfixed(-0.5968,1,L_SIZE),
				to_sfixed(-0.5965,1,L_SIZE),
				to_sfixed(-0.5963,1,L_SIZE),
				to_sfixed(-0.5961,1,L_SIZE),
				to_sfixed(-0.5958,1,L_SIZE),
				to_sfixed(-0.5956,1,L_SIZE),
				to_sfixed(-0.5954,1,L_SIZE),
				to_sfixed(-0.5951,1,L_SIZE),
				to_sfixed(-0.5949,1,L_SIZE),
				to_sfixed(-0.5946,1,L_SIZE),
				to_sfixed(-0.5944,1,L_SIZE),
				to_sfixed(-0.5942,1,L_SIZE),
				to_sfixed(-0.5939,1,L_SIZE),
				to_sfixed(-0.5937,1,L_SIZE),
				to_sfixed(-0.5935,1,L_SIZE),
				to_sfixed(-0.5932,1,L_SIZE),
				to_sfixed(-0.5930,1,L_SIZE),
				to_sfixed(-0.5927,1,L_SIZE),
				to_sfixed(-0.5925,1,L_SIZE),
				to_sfixed(-0.5923,1,L_SIZE),
				to_sfixed(-0.5920,1,L_SIZE),
				to_sfixed(-0.5918,1,L_SIZE),
				to_sfixed(-0.5916,1,L_SIZE),
				to_sfixed(-0.5913,1,L_SIZE),
				to_sfixed(-0.5911,1,L_SIZE),
				to_sfixed(-0.5908,1,L_SIZE),
				to_sfixed(-0.5906,1,L_SIZE),
				to_sfixed(-0.5904,1,L_SIZE),
				to_sfixed(-0.5901,1,L_SIZE),
				to_sfixed(-0.5899,1,L_SIZE),
				to_sfixed(-0.5896,1,L_SIZE),
				to_sfixed(-0.5894,1,L_SIZE),
				to_sfixed(-0.5892,1,L_SIZE),
				to_sfixed(-0.5889,1,L_SIZE),
				to_sfixed(-0.5887,1,L_SIZE),
				to_sfixed(-0.5885,1,L_SIZE),
				to_sfixed(-0.5882,1,L_SIZE),
				to_sfixed(-0.5880,1,L_SIZE),
				to_sfixed(-0.5877,1,L_SIZE),
				to_sfixed(-0.5875,1,L_SIZE),
				to_sfixed(-0.5873,1,L_SIZE),
				to_sfixed(-0.5870,1,L_SIZE),
				to_sfixed(-0.5868,1,L_SIZE),
				to_sfixed(-0.5865,1,L_SIZE),
				to_sfixed(-0.5863,1,L_SIZE),
				to_sfixed(-0.5861,1,L_SIZE),
				to_sfixed(-0.5858,1,L_SIZE),
				to_sfixed(-0.5856,1,L_SIZE),
				to_sfixed(-0.5853,1,L_SIZE),
				to_sfixed(-0.5851,1,L_SIZE),
				to_sfixed(-0.5848,1,L_SIZE),
				to_sfixed(-0.5846,1,L_SIZE),
				to_sfixed(-0.5844,1,L_SIZE),
				to_sfixed(-0.5841,1,L_SIZE),
				to_sfixed(-0.5839,1,L_SIZE),
				to_sfixed(-0.5836,1,L_SIZE),
				to_sfixed(-0.5834,1,L_SIZE),
				to_sfixed(-0.5832,1,L_SIZE),
				to_sfixed(-0.5829,1,L_SIZE),
				to_sfixed(-0.5827,1,L_SIZE),
				to_sfixed(-0.5824,1,L_SIZE),
				to_sfixed(-0.5822,1,L_SIZE),
				to_sfixed(-0.5819,1,L_SIZE),
				to_sfixed(-0.5817,1,L_SIZE),
				to_sfixed(-0.5815,1,L_SIZE),
				to_sfixed(-0.5812,1,L_SIZE),
				to_sfixed(-0.5810,1,L_SIZE),
				to_sfixed(-0.5807,1,L_SIZE),
				to_sfixed(-0.5805,1,L_SIZE),
				to_sfixed(-0.5803,1,L_SIZE),
				to_sfixed(-0.5800,1,L_SIZE),
				to_sfixed(-0.5798,1,L_SIZE),
				to_sfixed(-0.5795,1,L_SIZE),
				to_sfixed(-0.5793,1,L_SIZE),
				to_sfixed(-0.5790,1,L_SIZE),
				to_sfixed(-0.5788,1,L_SIZE),
				to_sfixed(-0.5785,1,L_SIZE),
				to_sfixed(-0.5783,1,L_SIZE),
				to_sfixed(-0.5781,1,L_SIZE),
				to_sfixed(-0.5778,1,L_SIZE),
				to_sfixed(-0.5776,1,L_SIZE),
				to_sfixed(-0.5773,1,L_SIZE),
				to_sfixed(-0.5771,1,L_SIZE),
				to_sfixed(-0.5768,1,L_SIZE),
				to_sfixed(-0.5766,1,L_SIZE),
				to_sfixed(-0.5764,1,L_SIZE),
				to_sfixed(-0.5761,1,L_SIZE),
				to_sfixed(-0.5759,1,L_SIZE),
				to_sfixed(-0.5756,1,L_SIZE),
				to_sfixed(-0.5754,1,L_SIZE),
				to_sfixed(-0.5751,1,L_SIZE),
				to_sfixed(-0.5749,1,L_SIZE),
				to_sfixed(-0.5746,1,L_SIZE),
				to_sfixed(-0.5744,1,L_SIZE),
				to_sfixed(-0.5741,1,L_SIZE),
				to_sfixed(-0.5739,1,L_SIZE),
				to_sfixed(-0.5737,1,L_SIZE),
				to_sfixed(-0.5734,1,L_SIZE),
				to_sfixed(-0.5732,1,L_SIZE),
				to_sfixed(-0.5729,1,L_SIZE),
				to_sfixed(-0.5727,1,L_SIZE),
				to_sfixed(-0.5724,1,L_SIZE),
				to_sfixed(-0.5722,1,L_SIZE),
				to_sfixed(-0.5719,1,L_SIZE),
				to_sfixed(-0.5717,1,L_SIZE),
				to_sfixed(-0.5714,1,L_SIZE),
				to_sfixed(-0.5712,1,L_SIZE),
				to_sfixed(-0.5709,1,L_SIZE),
				to_sfixed(-0.5707,1,L_SIZE),
				to_sfixed(-0.5705,1,L_SIZE),
				to_sfixed(-0.5702,1,L_SIZE),
				to_sfixed(-0.5700,1,L_SIZE),
				to_sfixed(-0.5697,1,L_SIZE),
				to_sfixed(-0.5695,1,L_SIZE),
				to_sfixed(-0.5692,1,L_SIZE),
				to_sfixed(-0.5690,1,L_SIZE),
				to_sfixed(-0.5687,1,L_SIZE),
				to_sfixed(-0.5685,1,L_SIZE),
				to_sfixed(-0.5682,1,L_SIZE),
				to_sfixed(-0.5680,1,L_SIZE),
				to_sfixed(-0.5677,1,L_SIZE),
				to_sfixed(-0.5675,1,L_SIZE),
				to_sfixed(-0.5672,1,L_SIZE),
				to_sfixed(-0.5670,1,L_SIZE),
				to_sfixed(-0.5667,1,L_SIZE),
				to_sfixed(-0.5665,1,L_SIZE),
				to_sfixed(-0.5662,1,L_SIZE),
				to_sfixed(-0.5660,1,L_SIZE),
				to_sfixed(-0.5657,1,L_SIZE),
				to_sfixed(-0.5655,1,L_SIZE),
				to_sfixed(-0.5652,1,L_SIZE),
				to_sfixed(-0.5650,1,L_SIZE),
				to_sfixed(-0.5647,1,L_SIZE),
				to_sfixed(-0.5645,1,L_SIZE),
				to_sfixed(-0.5642,1,L_SIZE),
				to_sfixed(-0.5640,1,L_SIZE),
				to_sfixed(-0.5637,1,L_SIZE),
				to_sfixed(-0.5635,1,L_SIZE),
				to_sfixed(-0.5632,1,L_SIZE),
				to_sfixed(-0.5630,1,L_SIZE),
				to_sfixed(-0.5627,1,L_SIZE),
				to_sfixed(-0.5625,1,L_SIZE),
				to_sfixed(-0.5622,1,L_SIZE),
				to_sfixed(-0.5620,1,L_SIZE),
				to_sfixed(-0.5617,1,L_SIZE),
				to_sfixed(-0.5615,1,L_SIZE),
				to_sfixed(-0.5612,1,L_SIZE),
				to_sfixed(-0.5610,1,L_SIZE),
				to_sfixed(-0.5607,1,L_SIZE),
				to_sfixed(-0.5605,1,L_SIZE),
				to_sfixed(-0.5602,1,L_SIZE),
				to_sfixed(-0.5600,1,L_SIZE),
				to_sfixed(-0.5597,1,L_SIZE),
				to_sfixed(-0.5595,1,L_SIZE),
				to_sfixed(-0.5592,1,L_SIZE),
				to_sfixed(-0.5590,1,L_SIZE),
				to_sfixed(-0.5587,1,L_SIZE),
				to_sfixed(-0.5585,1,L_SIZE),
				to_sfixed(-0.5582,1,L_SIZE),
				to_sfixed(-0.5580,1,L_SIZE),
				to_sfixed(-0.5577,1,L_SIZE),
				to_sfixed(-0.5575,1,L_SIZE),
				to_sfixed(-0.5572,1,L_SIZE),
				to_sfixed(-0.5570,1,L_SIZE),
				to_sfixed(-0.5567,1,L_SIZE),
				to_sfixed(-0.5565,1,L_SIZE),
				to_sfixed(-0.5562,1,L_SIZE),
				to_sfixed(-0.5560,1,L_SIZE),
				to_sfixed(-0.5557,1,L_SIZE),
				to_sfixed(-0.5554,1,L_SIZE),
				to_sfixed(-0.5552,1,L_SIZE),
				to_sfixed(-0.5549,1,L_SIZE),
				to_sfixed(-0.5547,1,L_SIZE),
				to_sfixed(-0.5544,1,L_SIZE),
				to_sfixed(-0.5542,1,L_SIZE),
				to_sfixed(-0.5539,1,L_SIZE),
				to_sfixed(-0.5537,1,L_SIZE),
				to_sfixed(-0.5534,1,L_SIZE),
				to_sfixed(-0.5532,1,L_SIZE),
				to_sfixed(-0.5529,1,L_SIZE),
				to_sfixed(-0.5527,1,L_SIZE),
				to_sfixed(-0.5524,1,L_SIZE),
				to_sfixed(-0.5521,1,L_SIZE),
				to_sfixed(-0.5519,1,L_SIZE),
				to_sfixed(-0.5516,1,L_SIZE),
				to_sfixed(-0.5514,1,L_SIZE),
				to_sfixed(-0.5511,1,L_SIZE),
				to_sfixed(-0.5509,1,L_SIZE),
				to_sfixed(-0.5506,1,L_SIZE),
				to_sfixed(-0.5504,1,L_SIZE),
				to_sfixed(-0.5501,1,L_SIZE),
				to_sfixed(-0.5498,1,L_SIZE),
				to_sfixed(-0.5496,1,L_SIZE),
				to_sfixed(-0.5493,1,L_SIZE),
				to_sfixed(-0.5491,1,L_SIZE),
				to_sfixed(-0.5488,1,L_SIZE),
				to_sfixed(-0.5486,1,L_SIZE),
				to_sfixed(-0.5483,1,L_SIZE),
				to_sfixed(-0.5481,1,L_SIZE),
				to_sfixed(-0.5478,1,L_SIZE),
				to_sfixed(-0.5475,1,L_SIZE),
				to_sfixed(-0.5473,1,L_SIZE),
				to_sfixed(-0.5470,1,L_SIZE),
				to_sfixed(-0.5468,1,L_SIZE),
				to_sfixed(-0.5465,1,L_SIZE),
				to_sfixed(-0.5463,1,L_SIZE),
				to_sfixed(-0.5460,1,L_SIZE),
				to_sfixed(-0.5457,1,L_SIZE),
				to_sfixed(-0.5455,1,L_SIZE),
				to_sfixed(-0.5452,1,L_SIZE),
				to_sfixed(-0.5450,1,L_SIZE),
				to_sfixed(-0.5447,1,L_SIZE),
				to_sfixed(-0.5445,1,L_SIZE),
				to_sfixed(-0.5442,1,L_SIZE),
				to_sfixed(-0.5439,1,L_SIZE),
				to_sfixed(-0.5437,1,L_SIZE),
				to_sfixed(-0.5434,1,L_SIZE),
				to_sfixed(-0.5432,1,L_SIZE),
				to_sfixed(-0.5429,1,L_SIZE),
				to_sfixed(-0.5427,1,L_SIZE),
				to_sfixed(-0.5424,1,L_SIZE),
				to_sfixed(-0.5421,1,L_SIZE),
				to_sfixed(-0.5419,1,L_SIZE),
				to_sfixed(-0.5416,1,L_SIZE),
				to_sfixed(-0.5414,1,L_SIZE),
				to_sfixed(-0.5411,1,L_SIZE),
				to_sfixed(-0.5408,1,L_SIZE),
				to_sfixed(-0.5406,1,L_SIZE),
				to_sfixed(-0.5403,1,L_SIZE),
				to_sfixed(-0.5401,1,L_SIZE),
				to_sfixed(-0.5398,1,L_SIZE),
				to_sfixed(-0.5395,1,L_SIZE),
				to_sfixed(-0.5393,1,L_SIZE),
				to_sfixed(-0.5390,1,L_SIZE),
				to_sfixed(-0.5388,1,L_SIZE),
				to_sfixed(-0.5385,1,L_SIZE),
				to_sfixed(-0.5382,1,L_SIZE),
				to_sfixed(-0.5380,1,L_SIZE),
				to_sfixed(-0.5377,1,L_SIZE),
				to_sfixed(-0.5375,1,L_SIZE),
				to_sfixed(-0.5372,1,L_SIZE),
				to_sfixed(-0.5369,1,L_SIZE),
				to_sfixed(-0.5367,1,L_SIZE),
				to_sfixed(-0.5364,1,L_SIZE),
				to_sfixed(-0.5362,1,L_SIZE),
				to_sfixed(-0.5359,1,L_SIZE),
				to_sfixed(-0.5356,1,L_SIZE),
				to_sfixed(-0.5354,1,L_SIZE),
				to_sfixed(-0.5351,1,L_SIZE),
				to_sfixed(-0.5349,1,L_SIZE),
				to_sfixed(-0.5346,1,L_SIZE),
				to_sfixed(-0.5343,1,L_SIZE),
				to_sfixed(-0.5341,1,L_SIZE),
				to_sfixed(-0.5338,1,L_SIZE),
				to_sfixed(-0.5335,1,L_SIZE),
				to_sfixed(-0.5333,1,L_SIZE),
				to_sfixed(-0.5330,1,L_SIZE),
				to_sfixed(-0.5328,1,L_SIZE),
				to_sfixed(-0.5325,1,L_SIZE),
				to_sfixed(-0.5322,1,L_SIZE),
				to_sfixed(-0.5320,1,L_SIZE),
				to_sfixed(-0.5317,1,L_SIZE),
				to_sfixed(-0.5314,1,L_SIZE),
				to_sfixed(-0.5312,1,L_SIZE),
				to_sfixed(-0.5309,1,L_SIZE),
				to_sfixed(-0.5307,1,L_SIZE),
				to_sfixed(-0.5304,1,L_SIZE),
				to_sfixed(-0.5301,1,L_SIZE),
				to_sfixed(-0.5299,1,L_SIZE),
				to_sfixed(-0.5296,1,L_SIZE),
				to_sfixed(-0.5293,1,L_SIZE),
				to_sfixed(-0.5291,1,L_SIZE),
				to_sfixed(-0.5288,1,L_SIZE),
				to_sfixed(-0.5286,1,L_SIZE),
				to_sfixed(-0.5283,1,L_SIZE),
				to_sfixed(-0.5280,1,L_SIZE),
				to_sfixed(-0.5278,1,L_SIZE),
				to_sfixed(-0.5275,1,L_SIZE),
				to_sfixed(-0.5272,1,L_SIZE),
				to_sfixed(-0.5270,1,L_SIZE),
				to_sfixed(-0.5267,1,L_SIZE),
				to_sfixed(-0.5264,1,L_SIZE),
				to_sfixed(-0.5262,1,L_SIZE),
				to_sfixed(-0.5259,1,L_SIZE),
				to_sfixed(-0.5256,1,L_SIZE),
				to_sfixed(-0.5254,1,L_SIZE),
				to_sfixed(-0.5251,1,L_SIZE),
				to_sfixed(-0.5248,1,L_SIZE),
				to_sfixed(-0.5246,1,L_SIZE),
				to_sfixed(-0.5243,1,L_SIZE),
				to_sfixed(-0.5241,1,L_SIZE),
				to_sfixed(-0.5238,1,L_SIZE),
				to_sfixed(-0.5235,1,L_SIZE),
				to_sfixed(-0.5233,1,L_SIZE),
				to_sfixed(-0.5230,1,L_SIZE),
				to_sfixed(-0.5227,1,L_SIZE),
				to_sfixed(-0.5225,1,L_SIZE),
				to_sfixed(-0.5222,1,L_SIZE),
				to_sfixed(-0.5219,1,L_SIZE),
				to_sfixed(-0.5217,1,L_SIZE),
				to_sfixed(-0.5214,1,L_SIZE),
				to_sfixed(-0.5211,1,L_SIZE),
				to_sfixed(-0.5209,1,L_SIZE),
				to_sfixed(-0.5206,1,L_SIZE),
				to_sfixed(-0.5203,1,L_SIZE),
				to_sfixed(-0.5201,1,L_SIZE),
				to_sfixed(-0.5198,1,L_SIZE),
				to_sfixed(-0.5195,1,L_SIZE),
				to_sfixed(-0.5193,1,L_SIZE),
				to_sfixed(-0.5190,1,L_SIZE),
				to_sfixed(-0.5187,1,L_SIZE),
				to_sfixed(-0.5185,1,L_SIZE),
				to_sfixed(-0.5182,1,L_SIZE),
				to_sfixed(-0.5179,1,L_SIZE),
				to_sfixed(-0.5176,1,L_SIZE),
				to_sfixed(-0.5174,1,L_SIZE),
				to_sfixed(-0.5171,1,L_SIZE),
				to_sfixed(-0.5168,1,L_SIZE),
				to_sfixed(-0.5166,1,L_SIZE),
				to_sfixed(-0.5163,1,L_SIZE),
				to_sfixed(-0.5160,1,L_SIZE),
				to_sfixed(-0.5158,1,L_SIZE),
				to_sfixed(-0.5155,1,L_SIZE),
				to_sfixed(-0.5152,1,L_SIZE),
				to_sfixed(-0.5150,1,L_SIZE),
				to_sfixed(-0.5147,1,L_SIZE),
				to_sfixed(-0.5144,1,L_SIZE),
				to_sfixed(-0.5142,1,L_SIZE),
				to_sfixed(-0.5139,1,L_SIZE),
				to_sfixed(-0.5136,1,L_SIZE),
				to_sfixed(-0.5133,1,L_SIZE),
				to_sfixed(-0.5131,1,L_SIZE),
				to_sfixed(-0.5128,1,L_SIZE),
				to_sfixed(-0.5125,1,L_SIZE),
				to_sfixed(-0.5123,1,L_SIZE),
				to_sfixed(-0.5120,1,L_SIZE),
				to_sfixed(-0.5117,1,L_SIZE),
				to_sfixed(-0.5115,1,L_SIZE),
				to_sfixed(-0.5112,1,L_SIZE),
				to_sfixed(-0.5109,1,L_SIZE),
				to_sfixed(-0.5106,1,L_SIZE),
				to_sfixed(-0.5104,1,L_SIZE),
				to_sfixed(-0.5101,1,L_SIZE),
				to_sfixed(-0.5098,1,L_SIZE),
				to_sfixed(-0.5096,1,L_SIZE),
				to_sfixed(-0.5093,1,L_SIZE),
				to_sfixed(-0.5090,1,L_SIZE),
				to_sfixed(-0.5087,1,L_SIZE),
				to_sfixed(-0.5085,1,L_SIZE),
				to_sfixed(-0.5082,1,L_SIZE),
				to_sfixed(-0.5079,1,L_SIZE),
				to_sfixed(-0.5077,1,L_SIZE),
				to_sfixed(-0.5074,1,L_SIZE),
				to_sfixed(-0.5071,1,L_SIZE),
				to_sfixed(-0.5068,1,L_SIZE),
				to_sfixed(-0.5066,1,L_SIZE),
				to_sfixed(-0.5063,1,L_SIZE),
				to_sfixed(-0.5060,1,L_SIZE),
				to_sfixed(-0.5058,1,L_SIZE),
				to_sfixed(-0.5055,1,L_SIZE),
				to_sfixed(-0.5052,1,L_SIZE),
				to_sfixed(-0.5049,1,L_SIZE),
				to_sfixed(-0.5047,1,L_SIZE),
				to_sfixed(-0.5044,1,L_SIZE),
				to_sfixed(-0.5041,1,L_SIZE),
				to_sfixed(-0.5038,1,L_SIZE),
				to_sfixed(-0.5036,1,L_SIZE),
				to_sfixed(-0.5033,1,L_SIZE),
				to_sfixed(-0.5030,1,L_SIZE),
				to_sfixed(-0.5027,1,L_SIZE),
				to_sfixed(-0.5025,1,L_SIZE),
				to_sfixed(-0.5022,1,L_SIZE),
				to_sfixed(-0.5019,1,L_SIZE),
				to_sfixed(-0.5017,1,L_SIZE),
				to_sfixed(-0.5014,1,L_SIZE),
				to_sfixed(-0.5011,1,L_SIZE),
				to_sfixed(-0.5008,1,L_SIZE),
				to_sfixed(-0.5006,1,L_SIZE),
				to_sfixed(-0.5003,1,L_SIZE),
				to_sfixed(-0.5000,1,L_SIZE),
				to_sfixed(-0.4997,1,L_SIZE),
				to_sfixed(-0.4995,1,L_SIZE),
				to_sfixed(-0.4992,1,L_SIZE),
				to_sfixed(-0.4989,1,L_SIZE),
				to_sfixed(-0.4986,1,L_SIZE),
				to_sfixed(-0.4984,1,L_SIZE),
				to_sfixed(-0.4981,1,L_SIZE),
				to_sfixed(-0.4978,1,L_SIZE),
				to_sfixed(-0.4975,1,L_SIZE),
				to_sfixed(-0.4973,1,L_SIZE),
				to_sfixed(-0.4970,1,L_SIZE),
				to_sfixed(-0.4967,1,L_SIZE),
				to_sfixed(-0.4964,1,L_SIZE),
				to_sfixed(-0.4962,1,L_SIZE),
				to_sfixed(-0.4959,1,L_SIZE),
				to_sfixed(-0.4956,1,L_SIZE),
				to_sfixed(-0.4953,1,L_SIZE),
				to_sfixed(-0.4950,1,L_SIZE),
				to_sfixed(-0.4948,1,L_SIZE),
				to_sfixed(-0.4945,1,L_SIZE),
				to_sfixed(-0.4942,1,L_SIZE),
				to_sfixed(-0.4939,1,L_SIZE),
				to_sfixed(-0.4937,1,L_SIZE),
				to_sfixed(-0.4934,1,L_SIZE),
				to_sfixed(-0.4931,1,L_SIZE),
				to_sfixed(-0.4928,1,L_SIZE),
				to_sfixed(-0.4926,1,L_SIZE),
				to_sfixed(-0.4923,1,L_SIZE),
				to_sfixed(-0.4920,1,L_SIZE),
				to_sfixed(-0.4917,1,L_SIZE),
				to_sfixed(-0.4914,1,L_SIZE),
				to_sfixed(-0.4912,1,L_SIZE),
				to_sfixed(-0.4909,1,L_SIZE),
				to_sfixed(-0.4906,1,L_SIZE),
				to_sfixed(-0.4903,1,L_SIZE),
				to_sfixed(-0.4901,1,L_SIZE),
				to_sfixed(-0.4898,1,L_SIZE),
				to_sfixed(-0.4895,1,L_SIZE),
				to_sfixed(-0.4892,1,L_SIZE),
				to_sfixed(-0.4889,1,L_SIZE),
				to_sfixed(-0.4887,1,L_SIZE),
				to_sfixed(-0.4884,1,L_SIZE),
				to_sfixed(-0.4881,1,L_SIZE),
				to_sfixed(-0.4878,1,L_SIZE),
				to_sfixed(-0.4875,1,L_SIZE),
				to_sfixed(-0.4873,1,L_SIZE),
				to_sfixed(-0.4870,1,L_SIZE),
				to_sfixed(-0.4867,1,L_SIZE),
				to_sfixed(-0.4864,1,L_SIZE),
				to_sfixed(-0.4861,1,L_SIZE),
				to_sfixed(-0.4859,1,L_SIZE),
				to_sfixed(-0.4856,1,L_SIZE),
				to_sfixed(-0.4853,1,L_SIZE),
				to_sfixed(-0.4850,1,L_SIZE),
				to_sfixed(-0.4848,1,L_SIZE),
				to_sfixed(-0.4845,1,L_SIZE),
				to_sfixed(-0.4842,1,L_SIZE),
				to_sfixed(-0.4839,1,L_SIZE),
				to_sfixed(-0.4836,1,L_SIZE),
				to_sfixed(-0.4833,1,L_SIZE),
				to_sfixed(-0.4831,1,L_SIZE),
				to_sfixed(-0.4828,1,L_SIZE),
				to_sfixed(-0.4825,1,L_SIZE),
				to_sfixed(-0.4822,1,L_SIZE),
				to_sfixed(-0.4819,1,L_SIZE),
				to_sfixed(-0.4817,1,L_SIZE),
				to_sfixed(-0.4814,1,L_SIZE),
				to_sfixed(-0.4811,1,L_SIZE),
				to_sfixed(-0.4808,1,L_SIZE),
				to_sfixed(-0.4805,1,L_SIZE),
				to_sfixed(-0.4803,1,L_SIZE),
				to_sfixed(-0.4800,1,L_SIZE),
				to_sfixed(-0.4797,1,L_SIZE),
				to_sfixed(-0.4794,1,L_SIZE),
				to_sfixed(-0.4791,1,L_SIZE),
				to_sfixed(-0.4788,1,L_SIZE),
				to_sfixed(-0.4786,1,L_SIZE),
				to_sfixed(-0.4783,1,L_SIZE),
				to_sfixed(-0.4780,1,L_SIZE),
				to_sfixed(-0.4777,1,L_SIZE),
				to_sfixed(-0.4774,1,L_SIZE),
				to_sfixed(-0.4771,1,L_SIZE),
				to_sfixed(-0.4769,1,L_SIZE),
				to_sfixed(-0.4766,1,L_SIZE),
				to_sfixed(-0.4763,1,L_SIZE),
				to_sfixed(-0.4760,1,L_SIZE),
				to_sfixed(-0.4757,1,L_SIZE),
				to_sfixed(-0.4755,1,L_SIZE),
				to_sfixed(-0.4752,1,L_SIZE),
				to_sfixed(-0.4749,1,L_SIZE),
				to_sfixed(-0.4746,1,L_SIZE),
				to_sfixed(-0.4743,1,L_SIZE),
				to_sfixed(-0.4740,1,L_SIZE),
				to_sfixed(-0.4737,1,L_SIZE),
				to_sfixed(-0.4735,1,L_SIZE),
				to_sfixed(-0.4732,1,L_SIZE),
				to_sfixed(-0.4729,1,L_SIZE),
				to_sfixed(-0.4726,1,L_SIZE),
				to_sfixed(-0.4723,1,L_SIZE),
				to_sfixed(-0.4720,1,L_SIZE),
				to_sfixed(-0.4718,1,L_SIZE),
				to_sfixed(-0.4715,1,L_SIZE),
				to_sfixed(-0.4712,1,L_SIZE),
				to_sfixed(-0.4709,1,L_SIZE),
				to_sfixed(-0.4706,1,L_SIZE),
				to_sfixed(-0.4703,1,L_SIZE),
				to_sfixed(-0.4700,1,L_SIZE),
				to_sfixed(-0.4698,1,L_SIZE),
				to_sfixed(-0.4695,1,L_SIZE),
				to_sfixed(-0.4692,1,L_SIZE),
				to_sfixed(-0.4689,1,L_SIZE),
				to_sfixed(-0.4686,1,L_SIZE),
				to_sfixed(-0.4683,1,L_SIZE),
				to_sfixed(-0.4680,1,L_SIZE),
				to_sfixed(-0.4678,1,L_SIZE),
				to_sfixed(-0.4675,1,L_SIZE),
				to_sfixed(-0.4672,1,L_SIZE),
				to_sfixed(-0.4669,1,L_SIZE),
				to_sfixed(-0.4666,1,L_SIZE),
				to_sfixed(-0.4663,1,L_SIZE),
				to_sfixed(-0.4660,1,L_SIZE),
				to_sfixed(-0.4658,1,L_SIZE),
				to_sfixed(-0.4655,1,L_SIZE),
				to_sfixed(-0.4652,1,L_SIZE),
				to_sfixed(-0.4649,1,L_SIZE),
				to_sfixed(-0.4646,1,L_SIZE),
				to_sfixed(-0.4643,1,L_SIZE),
				to_sfixed(-0.4640,1,L_SIZE),
				to_sfixed(-0.4637,1,L_SIZE),
				to_sfixed(-0.4635,1,L_SIZE),
				to_sfixed(-0.4632,1,L_SIZE),
				to_sfixed(-0.4629,1,L_SIZE),
				to_sfixed(-0.4626,1,L_SIZE),
				to_sfixed(-0.4623,1,L_SIZE),
				to_sfixed(-0.4620,1,L_SIZE),
				to_sfixed(-0.4617,1,L_SIZE),
				to_sfixed(-0.4614,1,L_SIZE),
				to_sfixed(-0.4612,1,L_SIZE),
				to_sfixed(-0.4609,1,L_SIZE),
				to_sfixed(-0.4606,1,L_SIZE),
				to_sfixed(-0.4603,1,L_SIZE),
				to_sfixed(-0.4600,1,L_SIZE),
				to_sfixed(-0.4597,1,L_SIZE),
				to_sfixed(-0.4594,1,L_SIZE),
				to_sfixed(-0.4591,1,L_SIZE),
				to_sfixed(-0.4588,1,L_SIZE),
				to_sfixed(-0.4586,1,L_SIZE),
				to_sfixed(-0.4583,1,L_SIZE),
				to_sfixed(-0.4580,1,L_SIZE),
				to_sfixed(-0.4577,1,L_SIZE),
				to_sfixed(-0.4574,1,L_SIZE),
				to_sfixed(-0.4571,1,L_SIZE),
				to_sfixed(-0.4568,1,L_SIZE),
				to_sfixed(-0.4565,1,L_SIZE),
				to_sfixed(-0.4562,1,L_SIZE),
				to_sfixed(-0.4560,1,L_SIZE),
				to_sfixed(-0.4557,1,L_SIZE),
				to_sfixed(-0.4554,1,L_SIZE),
				to_sfixed(-0.4551,1,L_SIZE),
				to_sfixed(-0.4548,1,L_SIZE),
				to_sfixed(-0.4545,1,L_SIZE),
				to_sfixed(-0.4542,1,L_SIZE),
				to_sfixed(-0.4539,1,L_SIZE),
				to_sfixed(-0.4536,1,L_SIZE),
				to_sfixed(-0.4533,1,L_SIZE),
				to_sfixed(-0.4530,1,L_SIZE),
				to_sfixed(-0.4528,1,L_SIZE),
				to_sfixed(-0.4525,1,L_SIZE),
				to_sfixed(-0.4522,1,L_SIZE),
				to_sfixed(-0.4519,1,L_SIZE),
				to_sfixed(-0.4516,1,L_SIZE),
				to_sfixed(-0.4513,1,L_SIZE),
				to_sfixed(-0.4510,1,L_SIZE),
				to_sfixed(-0.4507,1,L_SIZE),
				to_sfixed(-0.4504,1,L_SIZE),
				to_sfixed(-0.4501,1,L_SIZE),
				to_sfixed(-0.4498,1,L_SIZE),
				to_sfixed(-0.4495,1,L_SIZE),
				to_sfixed(-0.4493,1,L_SIZE),
				to_sfixed(-0.4490,1,L_SIZE),
				to_sfixed(-0.4487,1,L_SIZE),
				to_sfixed(-0.4484,1,L_SIZE),
				to_sfixed(-0.4481,1,L_SIZE),
				to_sfixed(-0.4478,1,L_SIZE),
				to_sfixed(-0.4475,1,L_SIZE),
				to_sfixed(-0.4472,1,L_SIZE),
				to_sfixed(-0.4469,1,L_SIZE),
				to_sfixed(-0.4466,1,L_SIZE),
				to_sfixed(-0.4463,1,L_SIZE),
				to_sfixed(-0.4460,1,L_SIZE),
				to_sfixed(-0.4457,1,L_SIZE),
				to_sfixed(-0.4454,1,L_SIZE),
				to_sfixed(-0.4452,1,L_SIZE),
				to_sfixed(-0.4449,1,L_SIZE),
				to_sfixed(-0.4446,1,L_SIZE),
				to_sfixed(-0.4443,1,L_SIZE),
				to_sfixed(-0.4440,1,L_SIZE),
				to_sfixed(-0.4437,1,L_SIZE),
				to_sfixed(-0.4434,1,L_SIZE),
				to_sfixed(-0.4431,1,L_SIZE),
				to_sfixed(-0.4428,1,L_SIZE),
				to_sfixed(-0.4425,1,L_SIZE),
				to_sfixed(-0.4422,1,L_SIZE),
				to_sfixed(-0.4419,1,L_SIZE),
				to_sfixed(-0.4416,1,L_SIZE),
				to_sfixed(-0.4413,1,L_SIZE),
				to_sfixed(-0.4410,1,L_SIZE),
				to_sfixed(-0.4407,1,L_SIZE),
				to_sfixed(-0.4404,1,L_SIZE),
				to_sfixed(-0.4401,1,L_SIZE),
				to_sfixed(-0.4399,1,L_SIZE),
				to_sfixed(-0.4396,1,L_SIZE),
				to_sfixed(-0.4393,1,L_SIZE),
				to_sfixed(-0.4390,1,L_SIZE),
				to_sfixed(-0.4387,1,L_SIZE),
				to_sfixed(-0.4384,1,L_SIZE),
				to_sfixed(-0.4381,1,L_SIZE),
				to_sfixed(-0.4378,1,L_SIZE),
				to_sfixed(-0.4375,1,L_SIZE),
				to_sfixed(-0.4372,1,L_SIZE),
				to_sfixed(-0.4369,1,L_SIZE),
				to_sfixed(-0.4366,1,L_SIZE),
				to_sfixed(-0.4363,1,L_SIZE),
				to_sfixed(-0.4360,1,L_SIZE),
				to_sfixed(-0.4357,1,L_SIZE),
				to_sfixed(-0.4354,1,L_SIZE),
				to_sfixed(-0.4351,1,L_SIZE),
				to_sfixed(-0.4348,1,L_SIZE),
				to_sfixed(-0.4345,1,L_SIZE),
				to_sfixed(-0.4342,1,L_SIZE),
				to_sfixed(-0.4339,1,L_SIZE),
				to_sfixed(-0.4336,1,L_SIZE),
				to_sfixed(-0.4333,1,L_SIZE),
				to_sfixed(-0.4330,1,L_SIZE),
				to_sfixed(-0.4327,1,L_SIZE),
				to_sfixed(-0.4324,1,L_SIZE),
				to_sfixed(-0.4321,1,L_SIZE),
				to_sfixed(-0.4318,1,L_SIZE),
				to_sfixed(-0.4315,1,L_SIZE),
				to_sfixed(-0.4312,1,L_SIZE),
				to_sfixed(-0.4309,1,L_SIZE),
				to_sfixed(-0.4306,1,L_SIZE),
				to_sfixed(-0.4304,1,L_SIZE),
				to_sfixed(-0.4301,1,L_SIZE),
				to_sfixed(-0.4298,1,L_SIZE),
				to_sfixed(-0.4295,1,L_SIZE),
				to_sfixed(-0.4292,1,L_SIZE),
				to_sfixed(-0.4289,1,L_SIZE),
				to_sfixed(-0.4286,1,L_SIZE),
				to_sfixed(-0.4283,1,L_SIZE),
				to_sfixed(-0.4280,1,L_SIZE),
				to_sfixed(-0.4277,1,L_SIZE),
				to_sfixed(-0.4274,1,L_SIZE),
				to_sfixed(-0.4271,1,L_SIZE),
				to_sfixed(-0.4268,1,L_SIZE),
				to_sfixed(-0.4265,1,L_SIZE),
				to_sfixed(-0.4262,1,L_SIZE),
				to_sfixed(-0.4259,1,L_SIZE),
				to_sfixed(-0.4256,1,L_SIZE),
				to_sfixed(-0.4253,1,L_SIZE),
				to_sfixed(-0.4250,1,L_SIZE),
				to_sfixed(-0.4247,1,L_SIZE),
				to_sfixed(-0.4244,1,L_SIZE),
				to_sfixed(-0.4241,1,L_SIZE),
				to_sfixed(-0.4238,1,L_SIZE),
				to_sfixed(-0.4235,1,L_SIZE),
				to_sfixed(-0.4232,1,L_SIZE),
				to_sfixed(-0.4229,1,L_SIZE),
				to_sfixed(-0.4226,1,L_SIZE),
				to_sfixed(-0.4223,1,L_SIZE),
				to_sfixed(-0.4220,1,L_SIZE),
				to_sfixed(-0.4217,1,L_SIZE),
				to_sfixed(-0.4214,1,L_SIZE),
				to_sfixed(-0.4211,1,L_SIZE),
				to_sfixed(-0.4208,1,L_SIZE),
				to_sfixed(-0.4205,1,L_SIZE),
				to_sfixed(-0.4202,1,L_SIZE),
				to_sfixed(-0.4198,1,L_SIZE),
				to_sfixed(-0.4195,1,L_SIZE),
				to_sfixed(-0.4192,1,L_SIZE),
				to_sfixed(-0.4189,1,L_SIZE),
				to_sfixed(-0.4186,1,L_SIZE),
				to_sfixed(-0.4183,1,L_SIZE),
				to_sfixed(-0.4180,1,L_SIZE),
				to_sfixed(-0.4177,1,L_SIZE),
				to_sfixed(-0.4174,1,L_SIZE),
				to_sfixed(-0.4171,1,L_SIZE),
				to_sfixed(-0.4168,1,L_SIZE),
				to_sfixed(-0.4165,1,L_SIZE),
				to_sfixed(-0.4162,1,L_SIZE),
				to_sfixed(-0.4159,1,L_SIZE),
				to_sfixed(-0.4156,1,L_SIZE),
				to_sfixed(-0.4153,1,L_SIZE),
				to_sfixed(-0.4150,1,L_SIZE),
				to_sfixed(-0.4147,1,L_SIZE),
				to_sfixed(-0.4144,1,L_SIZE),
				to_sfixed(-0.4141,1,L_SIZE),
				to_sfixed(-0.4138,1,L_SIZE),
				to_sfixed(-0.4135,1,L_SIZE),
				to_sfixed(-0.4132,1,L_SIZE),
				to_sfixed(-0.4129,1,L_SIZE),
				to_sfixed(-0.4126,1,L_SIZE),
				to_sfixed(-0.4123,1,L_SIZE),
				to_sfixed(-0.4120,1,L_SIZE),
				to_sfixed(-0.4117,1,L_SIZE),
				to_sfixed(-0.4114,1,L_SIZE),
				to_sfixed(-0.4111,1,L_SIZE),
				to_sfixed(-0.4108,1,L_SIZE),
				to_sfixed(-0.4105,1,L_SIZE),
				to_sfixed(-0.4101,1,L_SIZE),
				to_sfixed(-0.4098,1,L_SIZE),
				to_sfixed(-0.4095,1,L_SIZE),
				to_sfixed(-0.4092,1,L_SIZE),
				to_sfixed(-0.4089,1,L_SIZE),
				to_sfixed(-0.4086,1,L_SIZE),
				to_sfixed(-0.4083,1,L_SIZE),
				to_sfixed(-0.4080,1,L_SIZE),
				to_sfixed(-0.4077,1,L_SIZE),
				to_sfixed(-0.4074,1,L_SIZE),
				to_sfixed(-0.4071,1,L_SIZE),
				to_sfixed(-0.4068,1,L_SIZE),
				to_sfixed(-0.4065,1,L_SIZE),
				to_sfixed(-0.4062,1,L_SIZE),
				to_sfixed(-0.4059,1,L_SIZE),
				to_sfixed(-0.4056,1,L_SIZE),
				to_sfixed(-0.4053,1,L_SIZE),
				to_sfixed(-0.4050,1,L_SIZE),
				to_sfixed(-0.4047,1,L_SIZE),
				to_sfixed(-0.4043,1,L_SIZE),
				to_sfixed(-0.4040,1,L_SIZE),
				to_sfixed(-0.4037,1,L_SIZE),
				to_sfixed(-0.4034,1,L_SIZE),
				to_sfixed(-0.4031,1,L_SIZE),
				to_sfixed(-0.4028,1,L_SIZE),
				to_sfixed(-0.4025,1,L_SIZE),
				to_sfixed(-0.4022,1,L_SIZE),
				to_sfixed(-0.4019,1,L_SIZE),
				to_sfixed(-0.4016,1,L_SIZE),
				to_sfixed(-0.4013,1,L_SIZE),
				to_sfixed(-0.4010,1,L_SIZE),
				to_sfixed(-0.4007,1,L_SIZE),
				to_sfixed(-0.4004,1,L_SIZE),
				to_sfixed(-0.4000,1,L_SIZE),
				to_sfixed(-0.3997,1,L_SIZE),
				to_sfixed(-0.3994,1,L_SIZE),
				to_sfixed(-0.3991,1,L_SIZE),
				to_sfixed(-0.3988,1,L_SIZE),
				to_sfixed(-0.3985,1,L_SIZE),
				to_sfixed(-0.3982,1,L_SIZE),
				to_sfixed(-0.3979,1,L_SIZE),
				to_sfixed(-0.3976,1,L_SIZE),
				to_sfixed(-0.3973,1,L_SIZE),
				to_sfixed(-0.3970,1,L_SIZE),
				to_sfixed(-0.3967,1,L_SIZE),
				to_sfixed(-0.3964,1,L_SIZE),
				to_sfixed(-0.3960,1,L_SIZE),
				to_sfixed(-0.3957,1,L_SIZE),
				to_sfixed(-0.3954,1,L_SIZE),
				to_sfixed(-0.3951,1,L_SIZE),
				to_sfixed(-0.3948,1,L_SIZE),
				to_sfixed(-0.3945,1,L_SIZE),
				to_sfixed(-0.3942,1,L_SIZE),
				to_sfixed(-0.3939,1,L_SIZE),
				to_sfixed(-0.3936,1,L_SIZE),
				to_sfixed(-0.3933,1,L_SIZE),
				to_sfixed(-0.3929,1,L_SIZE),
				to_sfixed(-0.3926,1,L_SIZE),
				to_sfixed(-0.3923,1,L_SIZE),
				to_sfixed(-0.3920,1,L_SIZE),
				to_sfixed(-0.3917,1,L_SIZE),
				to_sfixed(-0.3914,1,L_SIZE),
				to_sfixed(-0.3911,1,L_SIZE),
				to_sfixed(-0.3908,1,L_SIZE),
				to_sfixed(-0.3905,1,L_SIZE),
				to_sfixed(-0.3902,1,L_SIZE),
				to_sfixed(-0.3898,1,L_SIZE),
				to_sfixed(-0.3895,1,L_SIZE),
				to_sfixed(-0.3892,1,L_SIZE),
				to_sfixed(-0.3889,1,L_SIZE),
				to_sfixed(-0.3886,1,L_SIZE),
				to_sfixed(-0.3883,1,L_SIZE),
				to_sfixed(-0.3880,1,L_SIZE),
				to_sfixed(-0.3877,1,L_SIZE),
				to_sfixed(-0.3874,1,L_SIZE),
				to_sfixed(-0.3870,1,L_SIZE),
				to_sfixed(-0.3867,1,L_SIZE),
				to_sfixed(-0.3864,1,L_SIZE),
				to_sfixed(-0.3861,1,L_SIZE),
				to_sfixed(-0.3858,1,L_SIZE),
				to_sfixed(-0.3855,1,L_SIZE),
				to_sfixed(-0.3852,1,L_SIZE),
				to_sfixed(-0.3849,1,L_SIZE),
				to_sfixed(-0.3846,1,L_SIZE),
				to_sfixed(-0.3842,1,L_SIZE),
				to_sfixed(-0.3839,1,L_SIZE),
				to_sfixed(-0.3836,1,L_SIZE),
				to_sfixed(-0.3833,1,L_SIZE),
				to_sfixed(-0.3830,1,L_SIZE),
				to_sfixed(-0.3827,1,L_SIZE),
				to_sfixed(-0.3824,1,L_SIZE),
				to_sfixed(-0.3821,1,L_SIZE),
				to_sfixed(-0.3817,1,L_SIZE),
				to_sfixed(-0.3814,1,L_SIZE),
				to_sfixed(-0.3811,1,L_SIZE),
				to_sfixed(-0.3808,1,L_SIZE),
				to_sfixed(-0.3805,1,L_SIZE),
				to_sfixed(-0.3802,1,L_SIZE),
				to_sfixed(-0.3799,1,L_SIZE),
				to_sfixed(-0.3796,1,L_SIZE),
				to_sfixed(-0.3792,1,L_SIZE),
				to_sfixed(-0.3789,1,L_SIZE),
				to_sfixed(-0.3786,1,L_SIZE),
				to_sfixed(-0.3783,1,L_SIZE),
				to_sfixed(-0.3780,1,L_SIZE),
				to_sfixed(-0.3777,1,L_SIZE),
				to_sfixed(-0.3774,1,L_SIZE),
				to_sfixed(-0.3770,1,L_SIZE),
				to_sfixed(-0.3767,1,L_SIZE),
				to_sfixed(-0.3764,1,L_SIZE),
				to_sfixed(-0.3761,1,L_SIZE),
				to_sfixed(-0.3758,1,L_SIZE),
				to_sfixed(-0.3755,1,L_SIZE),
				to_sfixed(-0.3752,1,L_SIZE),
				to_sfixed(-0.3748,1,L_SIZE),
				to_sfixed(-0.3745,1,L_SIZE),
				to_sfixed(-0.3742,1,L_SIZE),
				to_sfixed(-0.3739,1,L_SIZE),
				to_sfixed(-0.3736,1,L_SIZE),
				to_sfixed(-0.3733,1,L_SIZE),
				to_sfixed(-0.3730,1,L_SIZE),
				to_sfixed(-0.3726,1,L_SIZE),
				to_sfixed(-0.3723,1,L_SIZE),
				to_sfixed(-0.3720,1,L_SIZE),
				to_sfixed(-0.3717,1,L_SIZE),
				to_sfixed(-0.3714,1,L_SIZE),
				to_sfixed(-0.3711,1,L_SIZE),
				to_sfixed(-0.3707,1,L_SIZE),
				to_sfixed(-0.3704,1,L_SIZE),
				to_sfixed(-0.3701,1,L_SIZE),
				to_sfixed(-0.3698,1,L_SIZE),
				to_sfixed(-0.3695,1,L_SIZE),
				to_sfixed(-0.3692,1,L_SIZE),
				to_sfixed(-0.3688,1,L_SIZE),
				to_sfixed(-0.3685,1,L_SIZE),
				to_sfixed(-0.3682,1,L_SIZE),
				to_sfixed(-0.3679,1,L_SIZE),
				to_sfixed(-0.3676,1,L_SIZE),
				to_sfixed(-0.3673,1,L_SIZE),
				to_sfixed(-0.3669,1,L_SIZE),
				to_sfixed(-0.3666,1,L_SIZE),
				to_sfixed(-0.3663,1,L_SIZE),
				to_sfixed(-0.3660,1,L_SIZE),
				to_sfixed(-0.3657,1,L_SIZE),
				to_sfixed(-0.3654,1,L_SIZE),
				to_sfixed(-0.3650,1,L_SIZE),
				to_sfixed(-0.3647,1,L_SIZE),
				to_sfixed(-0.3644,1,L_SIZE),
				to_sfixed(-0.3641,1,L_SIZE),
				to_sfixed(-0.3638,1,L_SIZE),
				to_sfixed(-0.3635,1,L_SIZE),
				to_sfixed(-0.3631,1,L_SIZE),
				to_sfixed(-0.3628,1,L_SIZE),
				to_sfixed(-0.3625,1,L_SIZE),
				to_sfixed(-0.3622,1,L_SIZE),
				to_sfixed(-0.3619,1,L_SIZE),
				to_sfixed(-0.3615,1,L_SIZE),
				to_sfixed(-0.3612,1,L_SIZE),
				to_sfixed(-0.3609,1,L_SIZE),
				to_sfixed(-0.3606,1,L_SIZE),
				to_sfixed(-0.3603,1,L_SIZE),
				to_sfixed(-0.3600,1,L_SIZE),
				to_sfixed(-0.3596,1,L_SIZE),
				to_sfixed(-0.3593,1,L_SIZE),
				to_sfixed(-0.3590,1,L_SIZE),
				to_sfixed(-0.3587,1,L_SIZE),
				to_sfixed(-0.3584,1,L_SIZE),
				to_sfixed(-0.3580,1,L_SIZE),
				to_sfixed(-0.3577,1,L_SIZE),
				to_sfixed(-0.3574,1,L_SIZE),
				to_sfixed(-0.3571,1,L_SIZE),
				to_sfixed(-0.3568,1,L_SIZE),
				to_sfixed(-0.3564,1,L_SIZE),
				to_sfixed(-0.3561,1,L_SIZE),
				to_sfixed(-0.3558,1,L_SIZE),
				to_sfixed(-0.3555,1,L_SIZE),
				to_sfixed(-0.3552,1,L_SIZE),
				to_sfixed(-0.3548,1,L_SIZE),
				to_sfixed(-0.3545,1,L_SIZE),
				to_sfixed(-0.3542,1,L_SIZE),
				to_sfixed(-0.3539,1,L_SIZE),
				to_sfixed(-0.3536,1,L_SIZE),
				to_sfixed(-0.3532,1,L_SIZE),
				to_sfixed(-0.3529,1,L_SIZE),
				to_sfixed(-0.3526,1,L_SIZE),
				to_sfixed(-0.3523,1,L_SIZE),
				to_sfixed(-0.3520,1,L_SIZE),
				to_sfixed(-0.3516,1,L_SIZE),
				to_sfixed(-0.3513,1,L_SIZE),
				to_sfixed(-0.3510,1,L_SIZE),
				to_sfixed(-0.3507,1,L_SIZE),
				to_sfixed(-0.3504,1,L_SIZE),
				to_sfixed(-0.3500,1,L_SIZE),
				to_sfixed(-0.3497,1,L_SIZE),
				to_sfixed(-0.3494,1,L_SIZE),
				to_sfixed(-0.3491,1,L_SIZE),
				to_sfixed(-0.3487,1,L_SIZE),
				to_sfixed(-0.3484,1,L_SIZE),
				to_sfixed(-0.3481,1,L_SIZE),
				to_sfixed(-0.3478,1,L_SIZE),
				to_sfixed(-0.3475,1,L_SIZE),
				to_sfixed(-0.3471,1,L_SIZE),
				to_sfixed(-0.3468,1,L_SIZE),
				to_sfixed(-0.3465,1,L_SIZE),
				to_sfixed(-0.3462,1,L_SIZE),
				to_sfixed(-0.3458,1,L_SIZE),
				to_sfixed(-0.3455,1,L_SIZE),
				to_sfixed(-0.3452,1,L_SIZE),
				to_sfixed(-0.3449,1,L_SIZE),
				to_sfixed(-0.3446,1,L_SIZE),
				to_sfixed(-0.3442,1,L_SIZE),
				to_sfixed(-0.3439,1,L_SIZE),
				to_sfixed(-0.3436,1,L_SIZE),
				to_sfixed(-0.3433,1,L_SIZE),
				to_sfixed(-0.3429,1,L_SIZE),
				to_sfixed(-0.3426,1,L_SIZE),
				to_sfixed(-0.3423,1,L_SIZE),
				to_sfixed(-0.3420,1,L_SIZE),
				to_sfixed(-0.3416,1,L_SIZE),
				to_sfixed(-0.3413,1,L_SIZE),
				to_sfixed(-0.3410,1,L_SIZE),
				to_sfixed(-0.3407,1,L_SIZE),
				to_sfixed(-0.3404,1,L_SIZE),
				to_sfixed(-0.3400,1,L_SIZE),
				to_sfixed(-0.3397,1,L_SIZE),
				to_sfixed(-0.3394,1,L_SIZE),
				to_sfixed(-0.3391,1,L_SIZE),
				to_sfixed(-0.3387,1,L_SIZE),
				to_sfixed(-0.3384,1,L_SIZE),
				to_sfixed(-0.3381,1,L_SIZE),
				to_sfixed(-0.3378,1,L_SIZE),
				to_sfixed(-0.3374,1,L_SIZE),
				to_sfixed(-0.3371,1,L_SIZE),
				to_sfixed(-0.3368,1,L_SIZE),
				to_sfixed(-0.3365,1,L_SIZE),
				to_sfixed(-0.3361,1,L_SIZE),
				to_sfixed(-0.3358,1,L_SIZE),
				to_sfixed(-0.3355,1,L_SIZE),
				to_sfixed(-0.3352,1,L_SIZE),
				to_sfixed(-0.3348,1,L_SIZE),
				to_sfixed(-0.3345,1,L_SIZE),
				to_sfixed(-0.3342,1,L_SIZE),
				to_sfixed(-0.3339,1,L_SIZE),
				to_sfixed(-0.3335,1,L_SIZE),
				to_sfixed(-0.3332,1,L_SIZE),
				to_sfixed(-0.3329,1,L_SIZE),
				to_sfixed(-0.3326,1,L_SIZE),
				to_sfixed(-0.3322,1,L_SIZE),
				to_sfixed(-0.3319,1,L_SIZE),
				to_sfixed(-0.3316,1,L_SIZE),
				to_sfixed(-0.3313,1,L_SIZE),
				to_sfixed(-0.3309,1,L_SIZE),
				to_sfixed(-0.3306,1,L_SIZE),
				to_sfixed(-0.3303,1,L_SIZE),
				to_sfixed(-0.3300,1,L_SIZE),
				to_sfixed(-0.3296,1,L_SIZE),
				to_sfixed(-0.3293,1,L_SIZE),
				to_sfixed(-0.3290,1,L_SIZE),
				to_sfixed(-0.3286,1,L_SIZE),
				to_sfixed(-0.3283,1,L_SIZE),
				to_sfixed(-0.3280,1,L_SIZE),
				to_sfixed(-0.3277,1,L_SIZE),
				to_sfixed(-0.3273,1,L_SIZE),
				to_sfixed(-0.3270,1,L_SIZE),
				to_sfixed(-0.3267,1,L_SIZE),
				to_sfixed(-0.3264,1,L_SIZE),
				to_sfixed(-0.3260,1,L_SIZE),
				to_sfixed(-0.3257,1,L_SIZE),
				to_sfixed(-0.3254,1,L_SIZE),
				to_sfixed(-0.3250,1,L_SIZE),
				to_sfixed(-0.3247,1,L_SIZE),
				to_sfixed(-0.3244,1,L_SIZE),
				to_sfixed(-0.3241,1,L_SIZE),
				to_sfixed(-0.3237,1,L_SIZE),
				to_sfixed(-0.3234,1,L_SIZE),
				to_sfixed(-0.3231,1,L_SIZE),
				to_sfixed(-0.3228,1,L_SIZE),
				to_sfixed(-0.3224,1,L_SIZE),
				to_sfixed(-0.3221,1,L_SIZE),
				to_sfixed(-0.3218,1,L_SIZE),
				to_sfixed(-0.3214,1,L_SIZE),
				to_sfixed(-0.3211,1,L_SIZE),
				to_sfixed(-0.3208,1,L_SIZE),
				to_sfixed(-0.3205,1,L_SIZE),
				to_sfixed(-0.3201,1,L_SIZE),
				to_sfixed(-0.3198,1,L_SIZE),
				to_sfixed(-0.3195,1,L_SIZE),
				to_sfixed(-0.3191,1,L_SIZE),
				to_sfixed(-0.3188,1,L_SIZE),
				to_sfixed(-0.3185,1,L_SIZE),
				to_sfixed(-0.3182,1,L_SIZE),
				to_sfixed(-0.3178,1,L_SIZE),
				to_sfixed(-0.3175,1,L_SIZE),
				to_sfixed(-0.3172,1,L_SIZE),
				to_sfixed(-0.3168,1,L_SIZE),
				to_sfixed(-0.3165,1,L_SIZE),
				to_sfixed(-0.3162,1,L_SIZE),
				to_sfixed(-0.3158,1,L_SIZE),
				to_sfixed(-0.3155,1,L_SIZE),
				to_sfixed(-0.3152,1,L_SIZE),
				to_sfixed(-0.3149,1,L_SIZE),
				to_sfixed(-0.3145,1,L_SIZE),
				to_sfixed(-0.3142,1,L_SIZE),
				to_sfixed(-0.3139,1,L_SIZE),
				to_sfixed(-0.3135,1,L_SIZE),
				to_sfixed(-0.3132,1,L_SIZE),
				to_sfixed(-0.3129,1,L_SIZE),
				to_sfixed(-0.3125,1,L_SIZE),
				to_sfixed(-0.3122,1,L_SIZE),
				to_sfixed(-0.3119,1,L_SIZE),
				to_sfixed(-0.3116,1,L_SIZE),
				to_sfixed(-0.3112,1,L_SIZE),
				to_sfixed(-0.3109,1,L_SIZE),
				to_sfixed(-0.3106,1,L_SIZE),
				to_sfixed(-0.3102,1,L_SIZE),
				to_sfixed(-0.3099,1,L_SIZE),
				to_sfixed(-0.3096,1,L_SIZE),
				to_sfixed(-0.3092,1,L_SIZE),
				to_sfixed(-0.3089,1,L_SIZE),
				to_sfixed(-0.3086,1,L_SIZE),
				to_sfixed(-0.3082,1,L_SIZE),
				to_sfixed(-0.3079,1,L_SIZE),
				to_sfixed(-0.3076,1,L_SIZE),
				to_sfixed(-0.3072,1,L_SIZE),
				to_sfixed(-0.3069,1,L_SIZE),
				to_sfixed(-0.3066,1,L_SIZE),
				to_sfixed(-0.3063,1,L_SIZE),
				to_sfixed(-0.3059,1,L_SIZE),
				to_sfixed(-0.3056,1,L_SIZE),
				to_sfixed(-0.3053,1,L_SIZE),
				to_sfixed(-0.3049,1,L_SIZE),
				to_sfixed(-0.3046,1,L_SIZE),
				to_sfixed(-0.3043,1,L_SIZE),
				to_sfixed(-0.3039,1,L_SIZE),
				to_sfixed(-0.3036,1,L_SIZE),
				to_sfixed(-0.3033,1,L_SIZE),
				to_sfixed(-0.3029,1,L_SIZE),
				to_sfixed(-0.3026,1,L_SIZE),
				to_sfixed(-0.3023,1,L_SIZE),
				to_sfixed(-0.3019,1,L_SIZE),
				to_sfixed(-0.3016,1,L_SIZE),
				to_sfixed(-0.3013,1,L_SIZE),
				to_sfixed(-0.3009,1,L_SIZE),
				to_sfixed(-0.3006,1,L_SIZE),
				to_sfixed(-0.3003,1,L_SIZE),
				to_sfixed(-0.2999,1,L_SIZE),
				to_sfixed(-0.2996,1,L_SIZE),
				to_sfixed(-0.2993,1,L_SIZE),
				to_sfixed(-0.2989,1,L_SIZE),
				to_sfixed(-0.2986,1,L_SIZE),
				to_sfixed(-0.2983,1,L_SIZE),
				to_sfixed(-0.2979,1,L_SIZE),
				to_sfixed(-0.2976,1,L_SIZE),
				to_sfixed(-0.2973,1,L_SIZE),
				to_sfixed(-0.2969,1,L_SIZE),
				to_sfixed(-0.2966,1,L_SIZE),
				to_sfixed(-0.2963,1,L_SIZE),
				to_sfixed(-0.2959,1,L_SIZE),
				to_sfixed(-0.2956,1,L_SIZE),
				to_sfixed(-0.2953,1,L_SIZE),
				to_sfixed(-0.2949,1,L_SIZE),
				to_sfixed(-0.2946,1,L_SIZE),
				to_sfixed(-0.2943,1,L_SIZE),
				to_sfixed(-0.2939,1,L_SIZE),
				to_sfixed(-0.2936,1,L_SIZE),
				to_sfixed(-0.2933,1,L_SIZE),
				to_sfixed(-0.2929,1,L_SIZE),
				to_sfixed(-0.2926,1,L_SIZE),
				to_sfixed(-0.2923,1,L_SIZE),
				to_sfixed(-0.2919,1,L_SIZE),
				to_sfixed(-0.2916,1,L_SIZE),
				to_sfixed(-0.2912,1,L_SIZE),
				to_sfixed(-0.2909,1,L_SIZE),
				to_sfixed(-0.2906,1,L_SIZE),
				to_sfixed(-0.2902,1,L_SIZE),
				to_sfixed(-0.2899,1,L_SIZE),
				to_sfixed(-0.2896,1,L_SIZE),
				to_sfixed(-0.2892,1,L_SIZE),
				to_sfixed(-0.2889,1,L_SIZE),
				to_sfixed(-0.2886,1,L_SIZE),
				to_sfixed(-0.2882,1,L_SIZE),
				to_sfixed(-0.2879,1,L_SIZE),
				to_sfixed(-0.2876,1,L_SIZE),
				to_sfixed(-0.2872,1,L_SIZE),
				to_sfixed(-0.2869,1,L_SIZE),
				to_sfixed(-0.2865,1,L_SIZE),
				to_sfixed(-0.2862,1,L_SIZE),
				to_sfixed(-0.2859,1,L_SIZE),
				to_sfixed(-0.2855,1,L_SIZE),
				to_sfixed(-0.2852,1,L_SIZE),
				to_sfixed(-0.2849,1,L_SIZE),
				to_sfixed(-0.2845,1,L_SIZE),
				to_sfixed(-0.2842,1,L_SIZE),
				to_sfixed(-0.2839,1,L_SIZE),
				to_sfixed(-0.2835,1,L_SIZE),
				to_sfixed(-0.2832,1,L_SIZE),
				to_sfixed(-0.2828,1,L_SIZE),
				to_sfixed(-0.2825,1,L_SIZE),
				to_sfixed(-0.2822,1,L_SIZE),
				to_sfixed(-0.2818,1,L_SIZE),
				to_sfixed(-0.2815,1,L_SIZE),
				to_sfixed(-0.2812,1,L_SIZE),
				to_sfixed(-0.2808,1,L_SIZE),
				to_sfixed(-0.2805,1,L_SIZE),
				to_sfixed(-0.2801,1,L_SIZE),
				to_sfixed(-0.2798,1,L_SIZE),
				to_sfixed(-0.2795,1,L_SIZE),
				to_sfixed(-0.2791,1,L_SIZE),
				to_sfixed(-0.2788,1,L_SIZE),
				to_sfixed(-0.2785,1,L_SIZE),
				to_sfixed(-0.2781,1,L_SIZE),
				to_sfixed(-0.2778,1,L_SIZE),
				to_sfixed(-0.2774,1,L_SIZE),
				to_sfixed(-0.2771,1,L_SIZE),
				to_sfixed(-0.2768,1,L_SIZE),
				to_sfixed(-0.2764,1,L_SIZE),
				to_sfixed(-0.2761,1,L_SIZE),
				to_sfixed(-0.2758,1,L_SIZE),
				to_sfixed(-0.2754,1,L_SIZE),
				to_sfixed(-0.2751,1,L_SIZE),
				to_sfixed(-0.2747,1,L_SIZE),
				to_sfixed(-0.2744,1,L_SIZE),
				to_sfixed(-0.2741,1,L_SIZE),
				to_sfixed(-0.2737,1,L_SIZE),
				to_sfixed(-0.2734,1,L_SIZE),
				to_sfixed(-0.2730,1,L_SIZE),
				to_sfixed(-0.2727,1,L_SIZE),
				to_sfixed(-0.2724,1,L_SIZE),
				to_sfixed(-0.2720,1,L_SIZE),
				to_sfixed(-0.2717,1,L_SIZE),
				to_sfixed(-0.2713,1,L_SIZE),
				to_sfixed(-0.2710,1,L_SIZE),
				to_sfixed(-0.2707,1,L_SIZE),
				to_sfixed(-0.2703,1,L_SIZE),
				to_sfixed(-0.2700,1,L_SIZE),
				to_sfixed(-0.2697,1,L_SIZE),
				to_sfixed(-0.2693,1,L_SIZE),
				to_sfixed(-0.2690,1,L_SIZE),
				to_sfixed(-0.2686,1,L_SIZE),
				to_sfixed(-0.2683,1,L_SIZE),
				to_sfixed(-0.2680,1,L_SIZE),
				to_sfixed(-0.2676,1,L_SIZE),
				to_sfixed(-0.2673,1,L_SIZE),
				to_sfixed(-0.2669,1,L_SIZE),
				to_sfixed(-0.2666,1,L_SIZE),
				to_sfixed(-0.2663,1,L_SIZE),
				to_sfixed(-0.2659,1,L_SIZE),
				to_sfixed(-0.2656,1,L_SIZE),
				to_sfixed(-0.2652,1,L_SIZE),
				to_sfixed(-0.2649,1,L_SIZE),
				to_sfixed(-0.2646,1,L_SIZE),
				to_sfixed(-0.2642,1,L_SIZE),
				to_sfixed(-0.2639,1,L_SIZE),
				to_sfixed(-0.2635,1,L_SIZE),
				to_sfixed(-0.2632,1,L_SIZE),
				to_sfixed(-0.2628,1,L_SIZE),
				to_sfixed(-0.2625,1,L_SIZE),
				to_sfixed(-0.2622,1,L_SIZE),
				to_sfixed(-0.2618,1,L_SIZE),
				to_sfixed(-0.2615,1,L_SIZE),
				to_sfixed(-0.2611,1,L_SIZE),
				to_sfixed(-0.2608,1,L_SIZE),
				to_sfixed(-0.2605,1,L_SIZE),
				to_sfixed(-0.2601,1,L_SIZE),
				to_sfixed(-0.2598,1,L_SIZE),
				to_sfixed(-0.2594,1,L_SIZE),
				to_sfixed(-0.2591,1,L_SIZE),
				to_sfixed(-0.2588,1,L_SIZE),
				to_sfixed(-0.2584,1,L_SIZE),
				to_sfixed(-0.2581,1,L_SIZE),
				to_sfixed(-0.2577,1,L_SIZE),
				to_sfixed(-0.2574,1,L_SIZE),
				to_sfixed(-0.2570,1,L_SIZE),
				to_sfixed(-0.2567,1,L_SIZE),
				to_sfixed(-0.2564,1,L_SIZE),
				to_sfixed(-0.2560,1,L_SIZE),
				to_sfixed(-0.2557,1,L_SIZE),
				to_sfixed(-0.2553,1,L_SIZE),
				to_sfixed(-0.2550,1,L_SIZE),
				to_sfixed(-0.2546,1,L_SIZE),
				to_sfixed(-0.2543,1,L_SIZE),
				to_sfixed(-0.2540,1,L_SIZE),
				to_sfixed(-0.2536,1,L_SIZE),
				to_sfixed(-0.2533,1,L_SIZE),
				to_sfixed(-0.2529,1,L_SIZE),
				to_sfixed(-0.2526,1,L_SIZE),
				to_sfixed(-0.2522,1,L_SIZE),
				to_sfixed(-0.2519,1,L_SIZE),
				to_sfixed(-0.2516,1,L_SIZE),
				to_sfixed(-0.2512,1,L_SIZE),
				to_sfixed(-0.2509,1,L_SIZE),
				to_sfixed(-0.2505,1,L_SIZE),
				to_sfixed(-0.2502,1,L_SIZE),
				to_sfixed(-0.2498,1,L_SIZE),
				to_sfixed(-0.2495,1,L_SIZE),
				to_sfixed(-0.2492,1,L_SIZE),
				to_sfixed(-0.2488,1,L_SIZE),
				to_sfixed(-0.2485,1,L_SIZE),
				to_sfixed(-0.2481,1,L_SIZE),
				to_sfixed(-0.2478,1,L_SIZE),
				to_sfixed(-0.2474,1,L_SIZE),
				to_sfixed(-0.2471,1,L_SIZE),
				to_sfixed(-0.2468,1,L_SIZE),
				to_sfixed(-0.2464,1,L_SIZE),
				to_sfixed(-0.2461,1,L_SIZE),
				to_sfixed(-0.2457,1,L_SIZE),
				to_sfixed(-0.2454,1,L_SIZE),
				to_sfixed(-0.2450,1,L_SIZE),
				to_sfixed(-0.2447,1,L_SIZE),
				to_sfixed(-0.2443,1,L_SIZE),
				to_sfixed(-0.2440,1,L_SIZE),
				to_sfixed(-0.2437,1,L_SIZE),
				to_sfixed(-0.2433,1,L_SIZE),
				to_sfixed(-0.2430,1,L_SIZE),
				to_sfixed(-0.2426,1,L_SIZE),
				to_sfixed(-0.2423,1,L_SIZE),
				to_sfixed(-0.2419,1,L_SIZE),
				to_sfixed(-0.2416,1,L_SIZE),
				to_sfixed(-0.2412,1,L_SIZE),
				to_sfixed(-0.2409,1,L_SIZE),
				to_sfixed(-0.2406,1,L_SIZE),
				to_sfixed(-0.2402,1,L_SIZE),
				to_sfixed(-0.2399,1,L_SIZE),
				to_sfixed(-0.2395,1,L_SIZE),
				to_sfixed(-0.2392,1,L_SIZE),
				to_sfixed(-0.2388,1,L_SIZE),
				to_sfixed(-0.2385,1,L_SIZE),
				to_sfixed(-0.2381,1,L_SIZE),
				to_sfixed(-0.2378,1,L_SIZE),
				to_sfixed(-0.2374,1,L_SIZE),
				to_sfixed(-0.2371,1,L_SIZE),
				to_sfixed(-0.2368,1,L_SIZE),
				to_sfixed(-0.2364,1,L_SIZE),
				to_sfixed(-0.2361,1,L_SIZE),
				to_sfixed(-0.2357,1,L_SIZE),
				to_sfixed(-0.2354,1,L_SIZE),
				to_sfixed(-0.2350,1,L_SIZE),
				to_sfixed(-0.2347,1,L_SIZE),
				to_sfixed(-0.2343,1,L_SIZE),
				to_sfixed(-0.2340,1,L_SIZE),
				to_sfixed(-0.2336,1,L_SIZE),
				to_sfixed(-0.2333,1,L_SIZE),
				to_sfixed(-0.2329,1,L_SIZE),
				to_sfixed(-0.2326,1,L_SIZE),
				to_sfixed(-0.2323,1,L_SIZE),
				to_sfixed(-0.2319,1,L_SIZE),
				to_sfixed(-0.2316,1,L_SIZE),
				to_sfixed(-0.2312,1,L_SIZE),
				to_sfixed(-0.2309,1,L_SIZE),
				to_sfixed(-0.2305,1,L_SIZE),
				to_sfixed(-0.2302,1,L_SIZE),
				to_sfixed(-0.2298,1,L_SIZE),
				to_sfixed(-0.2295,1,L_SIZE),
				to_sfixed(-0.2291,1,L_SIZE),
				to_sfixed(-0.2288,1,L_SIZE),
				to_sfixed(-0.2284,1,L_SIZE),
				to_sfixed(-0.2281,1,L_SIZE),
				to_sfixed(-0.2277,1,L_SIZE),
				to_sfixed(-0.2274,1,L_SIZE),
				to_sfixed(-0.2271,1,L_SIZE),
				to_sfixed(-0.2267,1,L_SIZE),
				to_sfixed(-0.2264,1,L_SIZE),
				to_sfixed(-0.2260,1,L_SIZE),
				to_sfixed(-0.2257,1,L_SIZE),
				to_sfixed(-0.2253,1,L_SIZE),
				to_sfixed(-0.2250,1,L_SIZE),
				to_sfixed(-0.2246,1,L_SIZE),
				to_sfixed(-0.2243,1,L_SIZE),
				to_sfixed(-0.2239,1,L_SIZE),
				to_sfixed(-0.2236,1,L_SIZE),
				to_sfixed(-0.2232,1,L_SIZE),
				to_sfixed(-0.2229,1,L_SIZE),
				to_sfixed(-0.2225,1,L_SIZE),
				to_sfixed(-0.2222,1,L_SIZE),
				to_sfixed(-0.2218,1,L_SIZE),
				to_sfixed(-0.2215,1,L_SIZE),
				to_sfixed(-0.2211,1,L_SIZE),
				to_sfixed(-0.2208,1,L_SIZE),
				to_sfixed(-0.2204,1,L_SIZE),
				to_sfixed(-0.2201,1,L_SIZE),
				to_sfixed(-0.2197,1,L_SIZE),
				to_sfixed(-0.2194,1,L_SIZE),
				to_sfixed(-0.2190,1,L_SIZE),
				to_sfixed(-0.2187,1,L_SIZE),
				to_sfixed(-0.2184,1,L_SIZE),
				to_sfixed(-0.2180,1,L_SIZE),
				to_sfixed(-0.2177,1,L_SIZE),
				to_sfixed(-0.2173,1,L_SIZE),
				to_sfixed(-0.2170,1,L_SIZE),
				to_sfixed(-0.2166,1,L_SIZE),
				to_sfixed(-0.2163,1,L_SIZE),
				to_sfixed(-0.2159,1,L_SIZE),
				to_sfixed(-0.2156,1,L_SIZE),
				to_sfixed(-0.2152,1,L_SIZE),
				to_sfixed(-0.2149,1,L_SIZE),
				to_sfixed(-0.2145,1,L_SIZE),
				to_sfixed(-0.2142,1,L_SIZE),
				to_sfixed(-0.2138,1,L_SIZE),
				to_sfixed(-0.2135,1,L_SIZE),
				to_sfixed(-0.2131,1,L_SIZE),
				to_sfixed(-0.2128,1,L_SIZE),
				to_sfixed(-0.2124,1,L_SIZE),
				to_sfixed(-0.2121,1,L_SIZE),
				to_sfixed(-0.2117,1,L_SIZE),
				to_sfixed(-0.2114,1,L_SIZE),
				to_sfixed(-0.2110,1,L_SIZE),
				to_sfixed(-0.2107,1,L_SIZE),
				to_sfixed(-0.2103,1,L_SIZE),
				to_sfixed(-0.2100,1,L_SIZE),
				to_sfixed(-0.2096,1,L_SIZE),
				to_sfixed(-0.2093,1,L_SIZE),
				to_sfixed(-0.2089,1,L_SIZE),
				to_sfixed(-0.2086,1,L_SIZE),
				to_sfixed(-0.2082,1,L_SIZE),
				to_sfixed(-0.2079,1,L_SIZE),
				to_sfixed(-0.2075,1,L_SIZE),
				to_sfixed(-0.2072,1,L_SIZE),
				to_sfixed(-0.2068,1,L_SIZE),
				to_sfixed(-0.2065,1,L_SIZE),
				to_sfixed(-0.2061,1,L_SIZE),
				to_sfixed(-0.2058,1,L_SIZE),
				to_sfixed(-0.2054,1,L_SIZE),
				to_sfixed(-0.2051,1,L_SIZE),
				to_sfixed(-0.2047,1,L_SIZE),
				to_sfixed(-0.2044,1,L_SIZE),
				to_sfixed(-0.2040,1,L_SIZE),
				to_sfixed(-0.2037,1,L_SIZE),
				to_sfixed(-0.2033,1,L_SIZE),
				to_sfixed(-0.2030,1,L_SIZE),
				to_sfixed(-0.2026,1,L_SIZE),
				to_sfixed(-0.2023,1,L_SIZE),
				to_sfixed(-0.2019,1,L_SIZE),
				to_sfixed(-0.2015,1,L_SIZE),
				to_sfixed(-0.2012,1,L_SIZE),
				to_sfixed(-0.2008,1,L_SIZE),
				to_sfixed(-0.2005,1,L_SIZE),
				to_sfixed(-0.2001,1,L_SIZE),
				to_sfixed(-0.1998,1,L_SIZE),
				to_sfixed(-0.1994,1,L_SIZE),
				to_sfixed(-0.1991,1,L_SIZE),
				to_sfixed(-0.1987,1,L_SIZE),
				to_sfixed(-0.1984,1,L_SIZE),
				to_sfixed(-0.1980,1,L_SIZE),
				to_sfixed(-0.1977,1,L_SIZE),
				to_sfixed(-0.1973,1,L_SIZE),
				to_sfixed(-0.1970,1,L_SIZE),
				to_sfixed(-0.1966,1,L_SIZE),
				to_sfixed(-0.1963,1,L_SIZE),
				to_sfixed(-0.1959,1,L_SIZE),
				to_sfixed(-0.1956,1,L_SIZE),
				to_sfixed(-0.1952,1,L_SIZE),
				to_sfixed(-0.1949,1,L_SIZE),
				to_sfixed(-0.1945,1,L_SIZE),
				to_sfixed(-0.1942,1,L_SIZE),
				to_sfixed(-0.1938,1,L_SIZE),
				to_sfixed(-0.1935,1,L_SIZE),
				to_sfixed(-0.1931,1,L_SIZE),
				to_sfixed(-0.1927,1,L_SIZE),
				to_sfixed(-0.1924,1,L_SIZE),
				to_sfixed(-0.1920,1,L_SIZE),
				to_sfixed(-0.1917,1,L_SIZE),
				to_sfixed(-0.1913,1,L_SIZE),
				to_sfixed(-0.1910,1,L_SIZE),
				to_sfixed(-0.1906,1,L_SIZE),
				to_sfixed(-0.1903,1,L_SIZE),
				to_sfixed(-0.1899,1,L_SIZE),
				to_sfixed(-0.1896,1,L_SIZE),
				to_sfixed(-0.1892,1,L_SIZE),
				to_sfixed(-0.1889,1,L_SIZE),
				to_sfixed(-0.1885,1,L_SIZE),
				to_sfixed(-0.1882,1,L_SIZE),
				to_sfixed(-0.1878,1,L_SIZE),
				to_sfixed(-0.1875,1,L_SIZE),
				to_sfixed(-0.1871,1,L_SIZE),
				to_sfixed(-0.1867,1,L_SIZE),
				to_sfixed(-0.1864,1,L_SIZE),
				to_sfixed(-0.1860,1,L_SIZE),
				to_sfixed(-0.1857,1,L_SIZE),
				to_sfixed(-0.1853,1,L_SIZE),
				to_sfixed(-0.1850,1,L_SIZE),
				to_sfixed(-0.1846,1,L_SIZE),
				to_sfixed(-0.1843,1,L_SIZE),
				to_sfixed(-0.1839,1,L_SIZE),
				to_sfixed(-0.1836,1,L_SIZE),
				to_sfixed(-0.1832,1,L_SIZE),
				to_sfixed(-0.1829,1,L_SIZE),
				to_sfixed(-0.1825,1,L_SIZE),
				to_sfixed(-0.1821,1,L_SIZE),
				to_sfixed(-0.1818,1,L_SIZE),
				to_sfixed(-0.1814,1,L_SIZE),
				to_sfixed(-0.1811,1,L_SIZE),
				to_sfixed(-0.1807,1,L_SIZE),
				to_sfixed(-0.1804,1,L_SIZE),
				to_sfixed(-0.1800,1,L_SIZE),
				to_sfixed(-0.1797,1,L_SIZE),
				to_sfixed(-0.1793,1,L_SIZE),
				to_sfixed(-0.1790,1,L_SIZE),
				to_sfixed(-0.1786,1,L_SIZE),
				to_sfixed(-0.1783,1,L_SIZE),
				to_sfixed(-0.1779,1,L_SIZE),
				to_sfixed(-0.1775,1,L_SIZE),
				to_sfixed(-0.1772,1,L_SIZE),
				to_sfixed(-0.1768,1,L_SIZE),
				to_sfixed(-0.1765,1,L_SIZE),
				to_sfixed(-0.1761,1,L_SIZE),
				to_sfixed(-0.1758,1,L_SIZE),
				to_sfixed(-0.1754,1,L_SIZE),
				to_sfixed(-0.1751,1,L_SIZE),
				to_sfixed(-0.1747,1,L_SIZE),
				to_sfixed(-0.1743,1,L_SIZE),
				to_sfixed(-0.1740,1,L_SIZE),
				to_sfixed(-0.1736,1,L_SIZE),
				to_sfixed(-0.1733,1,L_SIZE),
				to_sfixed(-0.1729,1,L_SIZE),
				to_sfixed(-0.1726,1,L_SIZE),
				to_sfixed(-0.1722,1,L_SIZE),
				to_sfixed(-0.1719,1,L_SIZE),
				to_sfixed(-0.1715,1,L_SIZE),
				to_sfixed(-0.1712,1,L_SIZE),
				to_sfixed(-0.1708,1,L_SIZE),
				to_sfixed(-0.1704,1,L_SIZE),
				to_sfixed(-0.1701,1,L_SIZE),
				to_sfixed(-0.1697,1,L_SIZE),
				to_sfixed(-0.1694,1,L_SIZE),
				to_sfixed(-0.1690,1,L_SIZE),
				to_sfixed(-0.1687,1,L_SIZE),
				to_sfixed(-0.1683,1,L_SIZE),
				to_sfixed(-0.1679,1,L_SIZE),
				to_sfixed(-0.1676,1,L_SIZE),
				to_sfixed(-0.1672,1,L_SIZE),
				to_sfixed(-0.1669,1,L_SIZE),
				to_sfixed(-0.1665,1,L_SIZE),
				to_sfixed(-0.1662,1,L_SIZE),
				to_sfixed(-0.1658,1,L_SIZE),
				to_sfixed(-0.1655,1,L_SIZE),
				to_sfixed(-0.1651,1,L_SIZE),
				to_sfixed(-0.1647,1,L_SIZE),
				to_sfixed(-0.1644,1,L_SIZE),
				to_sfixed(-0.1640,1,L_SIZE),
				to_sfixed(-0.1637,1,L_SIZE),
				to_sfixed(-0.1633,1,L_SIZE),
				to_sfixed(-0.1630,1,L_SIZE),
				to_sfixed(-0.1626,1,L_SIZE),
				to_sfixed(-0.1622,1,L_SIZE),
				to_sfixed(-0.1619,1,L_SIZE),
				to_sfixed(-0.1615,1,L_SIZE),
				to_sfixed(-0.1612,1,L_SIZE),
				to_sfixed(-0.1608,1,L_SIZE),
				to_sfixed(-0.1605,1,L_SIZE),
				to_sfixed(-0.1601,1,L_SIZE),
				to_sfixed(-0.1598,1,L_SIZE),
				to_sfixed(-0.1594,1,L_SIZE),
				to_sfixed(-0.1590,1,L_SIZE),
				to_sfixed(-0.1587,1,L_SIZE),
				to_sfixed(-0.1583,1,L_SIZE),
				to_sfixed(-0.1580,1,L_SIZE),
				to_sfixed(-0.1576,1,L_SIZE),
				to_sfixed(-0.1573,1,L_SIZE),
				to_sfixed(-0.1569,1,L_SIZE),
				to_sfixed(-0.1565,1,L_SIZE),
				to_sfixed(-0.1562,1,L_SIZE),
				to_sfixed(-0.1558,1,L_SIZE),
				to_sfixed(-0.1555,1,L_SIZE),
				to_sfixed(-0.1551,1,L_SIZE),
				to_sfixed(-0.1548,1,L_SIZE),
				to_sfixed(-0.1544,1,L_SIZE),
				to_sfixed(-0.1540,1,L_SIZE),
				to_sfixed(-0.1537,1,L_SIZE),
				to_sfixed(-0.1533,1,L_SIZE),
				to_sfixed(-0.1530,1,L_SIZE),
				to_sfixed(-0.1526,1,L_SIZE),
				to_sfixed(-0.1522,1,L_SIZE),
				to_sfixed(-0.1519,1,L_SIZE),
				to_sfixed(-0.1515,1,L_SIZE),
				to_sfixed(-0.1512,1,L_SIZE),
				to_sfixed(-0.1508,1,L_SIZE),
				to_sfixed(-0.1505,1,L_SIZE),
				to_sfixed(-0.1501,1,L_SIZE),
				to_sfixed(-0.1497,1,L_SIZE),
				to_sfixed(-0.1494,1,L_SIZE),
				to_sfixed(-0.1490,1,L_SIZE),
				to_sfixed(-0.1487,1,L_SIZE),
				to_sfixed(-0.1483,1,L_SIZE),
				to_sfixed(-0.1480,1,L_SIZE),
				to_sfixed(-0.1476,1,L_SIZE),
				to_sfixed(-0.1472,1,L_SIZE),
				to_sfixed(-0.1469,1,L_SIZE),
				to_sfixed(-0.1465,1,L_SIZE),
				to_sfixed(-0.1462,1,L_SIZE),
				to_sfixed(-0.1458,1,L_SIZE),
				to_sfixed(-0.1454,1,L_SIZE),
				to_sfixed(-0.1451,1,L_SIZE),
				to_sfixed(-0.1447,1,L_SIZE),
				to_sfixed(-0.1444,1,L_SIZE),
				to_sfixed(-0.1440,1,L_SIZE),
				to_sfixed(-0.1437,1,L_SIZE),
				to_sfixed(-0.1433,1,L_SIZE),
				to_sfixed(-0.1429,1,L_SIZE),
				to_sfixed(-0.1426,1,L_SIZE),
				to_sfixed(-0.1422,1,L_SIZE),
				to_sfixed(-0.1419,1,L_SIZE),
				to_sfixed(-0.1415,1,L_SIZE),
				to_sfixed(-0.1411,1,L_SIZE),
				to_sfixed(-0.1408,1,L_SIZE),
				to_sfixed(-0.1404,1,L_SIZE),
				to_sfixed(-0.1401,1,L_SIZE),
				to_sfixed(-0.1397,1,L_SIZE),
				to_sfixed(-0.1393,1,L_SIZE),
				to_sfixed(-0.1390,1,L_SIZE),
				to_sfixed(-0.1386,1,L_SIZE),
				to_sfixed(-0.1383,1,L_SIZE),
				to_sfixed(-0.1379,1,L_SIZE),
				to_sfixed(-0.1376,1,L_SIZE),
				to_sfixed(-0.1372,1,L_SIZE),
				to_sfixed(-0.1368,1,L_SIZE),
				to_sfixed(-0.1365,1,L_SIZE),
				to_sfixed(-0.1361,1,L_SIZE),
				to_sfixed(-0.1358,1,L_SIZE),
				to_sfixed(-0.1354,1,L_SIZE),
				to_sfixed(-0.1350,1,L_SIZE),
				to_sfixed(-0.1347,1,L_SIZE),
				to_sfixed(-0.1343,1,L_SIZE),
				to_sfixed(-0.1340,1,L_SIZE),
				to_sfixed(-0.1336,1,L_SIZE),
				to_sfixed(-0.1332,1,L_SIZE),
				to_sfixed(-0.1329,1,L_SIZE),
				to_sfixed(-0.1325,1,L_SIZE),
				to_sfixed(-0.1322,1,L_SIZE),
				to_sfixed(-0.1318,1,L_SIZE),
				to_sfixed(-0.1314,1,L_SIZE),
				to_sfixed(-0.1311,1,L_SIZE),
				to_sfixed(-0.1307,1,L_SIZE),
				to_sfixed(-0.1304,1,L_SIZE),
				to_sfixed(-0.1300,1,L_SIZE),
				to_sfixed(-0.1296,1,L_SIZE),
				to_sfixed(-0.1293,1,L_SIZE),
				to_sfixed(-0.1289,1,L_SIZE),
				to_sfixed(-0.1286,1,L_SIZE),
				to_sfixed(-0.1282,1,L_SIZE),
				to_sfixed(-0.1278,1,L_SIZE),
				to_sfixed(-0.1275,1,L_SIZE),
				to_sfixed(-0.1271,1,L_SIZE),
				to_sfixed(-0.1268,1,L_SIZE),
				to_sfixed(-0.1264,1,L_SIZE),
				to_sfixed(-0.1260,1,L_SIZE),
				to_sfixed(-0.1257,1,L_SIZE),
				to_sfixed(-0.1253,1,L_SIZE),
				to_sfixed(-0.1250,1,L_SIZE),
				to_sfixed(-0.1246,1,L_SIZE),
				to_sfixed(-0.1242,1,L_SIZE),
				to_sfixed(-0.1239,1,L_SIZE),
				to_sfixed(-0.1235,1,L_SIZE),
				to_sfixed(-0.1232,1,L_SIZE),
				to_sfixed(-0.1228,1,L_SIZE),
				to_sfixed(-0.1224,1,L_SIZE),
				to_sfixed(-0.1221,1,L_SIZE),
				to_sfixed(-0.1217,1,L_SIZE),
				to_sfixed(-0.1213,1,L_SIZE),
				to_sfixed(-0.1210,1,L_SIZE),
				to_sfixed(-0.1206,1,L_SIZE),
				to_sfixed(-0.1203,1,L_SIZE),
				to_sfixed(-0.1199,1,L_SIZE),
				to_sfixed(-0.1195,1,L_SIZE),
				to_sfixed(-0.1192,1,L_SIZE),
				to_sfixed(-0.1188,1,L_SIZE),
				to_sfixed(-0.1185,1,L_SIZE),
				to_sfixed(-0.1181,1,L_SIZE),
				to_sfixed(-0.1177,1,L_SIZE),
				to_sfixed(-0.1174,1,L_SIZE),
				to_sfixed(-0.1170,1,L_SIZE),
				to_sfixed(-0.1167,1,L_SIZE),
				to_sfixed(-0.1163,1,L_SIZE),
				to_sfixed(-0.1159,1,L_SIZE),
				to_sfixed(-0.1156,1,L_SIZE),
				to_sfixed(-0.1152,1,L_SIZE),
				to_sfixed(-0.1148,1,L_SIZE),
				to_sfixed(-0.1145,1,L_SIZE),
				to_sfixed(-0.1141,1,L_SIZE),
				to_sfixed(-0.1138,1,L_SIZE),
				to_sfixed(-0.1134,1,L_SIZE),
				to_sfixed(-0.1130,1,L_SIZE),
				to_sfixed(-0.1127,1,L_SIZE),
				to_sfixed(-0.1123,1,L_SIZE),
				to_sfixed(-0.1120,1,L_SIZE),
				to_sfixed(-0.1116,1,L_SIZE),
				to_sfixed(-0.1112,1,L_SIZE),
				to_sfixed(-0.1109,1,L_SIZE),
				to_sfixed(-0.1105,1,L_SIZE),
				to_sfixed(-0.1101,1,L_SIZE),
				to_sfixed(-0.1098,1,L_SIZE),
				to_sfixed(-0.1094,1,L_SIZE),
				to_sfixed(-0.1091,1,L_SIZE),
				to_sfixed(-0.1087,1,L_SIZE),
				to_sfixed(-0.1083,1,L_SIZE),
				to_sfixed(-0.1080,1,L_SIZE),
				to_sfixed(-0.1076,1,L_SIZE),
				to_sfixed(-0.1073,1,L_SIZE),
				to_sfixed(-0.1069,1,L_SIZE),
				to_sfixed(-0.1065,1,L_SIZE),
				to_sfixed(-0.1062,1,L_SIZE),
				to_sfixed(-0.1058,1,L_SIZE),
				to_sfixed(-0.1054,1,L_SIZE),
				to_sfixed(-0.1051,1,L_SIZE),
				to_sfixed(-0.1047,1,L_SIZE),
				to_sfixed(-0.1044,1,L_SIZE),
				to_sfixed(-0.1040,1,L_SIZE),
				to_sfixed(-0.1036,1,L_SIZE),
				to_sfixed(-0.1033,1,L_SIZE),
				to_sfixed(-0.1029,1,L_SIZE),
				to_sfixed(-0.1025,1,L_SIZE),
				to_sfixed(-0.1022,1,L_SIZE),
				to_sfixed(-0.1018,1,L_SIZE),
				to_sfixed(-0.1015,1,L_SIZE),
				to_sfixed(-0.1011,1,L_SIZE),
				to_sfixed(-0.1007,1,L_SIZE),
				to_sfixed(-0.1004,1,L_SIZE),
				to_sfixed(-0.1000,1,L_SIZE),
				to_sfixed(-0.0996,1,L_SIZE),
				to_sfixed(-0.0993,1,L_SIZE),
				to_sfixed(-0.0989,1,L_SIZE),
				to_sfixed(-0.0986,1,L_SIZE),
				to_sfixed(-0.0982,1,L_SIZE),
				to_sfixed(-0.0978,1,L_SIZE),
				to_sfixed(-0.0975,1,L_SIZE),
				to_sfixed(-0.0971,1,L_SIZE),
				to_sfixed(-0.0967,1,L_SIZE),
				to_sfixed(-0.0964,1,L_SIZE),
				to_sfixed(-0.0960,1,L_SIZE),
				to_sfixed(-0.0957,1,L_SIZE),
				to_sfixed(-0.0953,1,L_SIZE),
				to_sfixed(-0.0949,1,L_SIZE),
				to_sfixed(-0.0946,1,L_SIZE),
				to_sfixed(-0.0942,1,L_SIZE),
				to_sfixed(-0.0938,1,L_SIZE),
				to_sfixed(-0.0935,1,L_SIZE),
				to_sfixed(-0.0931,1,L_SIZE),
				to_sfixed(-0.0928,1,L_SIZE),
				to_sfixed(-0.0924,1,L_SIZE),
				to_sfixed(-0.0920,1,L_SIZE),
				to_sfixed(-0.0917,1,L_SIZE),
				to_sfixed(-0.0913,1,L_SIZE),
				to_sfixed(-0.0909,1,L_SIZE),
				to_sfixed(-0.0906,1,L_SIZE),
				to_sfixed(-0.0902,1,L_SIZE),
				to_sfixed(-0.0898,1,L_SIZE),
				to_sfixed(-0.0895,1,L_SIZE),
				to_sfixed(-0.0891,1,L_SIZE),
				to_sfixed(-0.0888,1,L_SIZE),
				to_sfixed(-0.0884,1,L_SIZE),
				to_sfixed(-0.0880,1,L_SIZE),
				to_sfixed(-0.0877,1,L_SIZE),
				to_sfixed(-0.0873,1,L_SIZE),
				to_sfixed(-0.0869,1,L_SIZE),
				to_sfixed(-0.0866,1,L_SIZE),
				to_sfixed(-0.0862,1,L_SIZE),
				to_sfixed(-0.0858,1,L_SIZE),
				to_sfixed(-0.0855,1,L_SIZE),
				to_sfixed(-0.0851,1,L_SIZE),
				to_sfixed(-0.0848,1,L_SIZE),
				to_sfixed(-0.0844,1,L_SIZE),
				to_sfixed(-0.0840,1,L_SIZE),
				to_sfixed(-0.0837,1,L_SIZE),
				to_sfixed(-0.0833,1,L_SIZE),
				to_sfixed(-0.0829,1,L_SIZE),
				to_sfixed(-0.0826,1,L_SIZE),
				to_sfixed(-0.0822,1,L_SIZE),
				to_sfixed(-0.0818,1,L_SIZE),
				to_sfixed(-0.0815,1,L_SIZE),
				to_sfixed(-0.0811,1,L_SIZE),
				to_sfixed(-0.0808,1,L_SIZE),
				to_sfixed(-0.0804,1,L_SIZE),
				to_sfixed(-0.0800,1,L_SIZE),
				to_sfixed(-0.0797,1,L_SIZE),
				to_sfixed(-0.0793,1,L_SIZE),
				to_sfixed(-0.0789,1,L_SIZE),
				to_sfixed(-0.0786,1,L_SIZE),
				to_sfixed(-0.0782,1,L_SIZE),
				to_sfixed(-0.0778,1,L_SIZE),
				to_sfixed(-0.0775,1,L_SIZE),
				to_sfixed(-0.0771,1,L_SIZE),
				to_sfixed(-0.0768,1,L_SIZE),
				to_sfixed(-0.0764,1,L_SIZE),
				to_sfixed(-0.0760,1,L_SIZE),
				to_sfixed(-0.0757,1,L_SIZE),
				to_sfixed(-0.0753,1,L_SIZE),
				to_sfixed(-0.0749,1,L_SIZE),
				to_sfixed(-0.0746,1,L_SIZE),
				to_sfixed(-0.0742,1,L_SIZE),
				to_sfixed(-0.0738,1,L_SIZE),
				to_sfixed(-0.0735,1,L_SIZE),
				to_sfixed(-0.0731,1,L_SIZE),
				to_sfixed(-0.0727,1,L_SIZE),
				to_sfixed(-0.0724,1,L_SIZE),
				to_sfixed(-0.0720,1,L_SIZE),
				to_sfixed(-0.0717,1,L_SIZE),
				to_sfixed(-0.0713,1,L_SIZE),
				to_sfixed(-0.0709,1,L_SIZE),
				to_sfixed(-0.0706,1,L_SIZE),
				to_sfixed(-0.0702,1,L_SIZE),
				to_sfixed(-0.0698,1,L_SIZE),
				to_sfixed(-0.0695,1,L_SIZE),
				to_sfixed(-0.0691,1,L_SIZE),
				to_sfixed(-0.0687,1,L_SIZE),
				to_sfixed(-0.0684,1,L_SIZE),
				to_sfixed(-0.0680,1,L_SIZE),
				to_sfixed(-0.0676,1,L_SIZE),
				to_sfixed(-0.0673,1,L_SIZE),
				to_sfixed(-0.0669,1,L_SIZE),
				to_sfixed(-0.0666,1,L_SIZE),
				to_sfixed(-0.0662,1,L_SIZE),
				to_sfixed(-0.0658,1,L_SIZE),
				to_sfixed(-0.0655,1,L_SIZE),
				to_sfixed(-0.0651,1,L_SIZE),
				to_sfixed(-0.0647,1,L_SIZE),
				to_sfixed(-0.0644,1,L_SIZE),
				to_sfixed(-0.0640,1,L_SIZE),
				to_sfixed(-0.0636,1,L_SIZE),
				to_sfixed(-0.0633,1,L_SIZE),
				to_sfixed(-0.0629,1,L_SIZE),
				to_sfixed(-0.0625,1,L_SIZE),
				to_sfixed(-0.0622,1,L_SIZE),
				to_sfixed(-0.0618,1,L_SIZE),
				to_sfixed(-0.0614,1,L_SIZE),
				to_sfixed(-0.0611,1,L_SIZE),
				to_sfixed(-0.0607,1,L_SIZE),
				to_sfixed(-0.0604,1,L_SIZE),
				to_sfixed(-0.0600,1,L_SIZE),
				to_sfixed(-0.0596,1,L_SIZE),
				to_sfixed(-0.0593,1,L_SIZE),
				to_sfixed(-0.0589,1,L_SIZE),
				to_sfixed(-0.0585,1,L_SIZE),
				to_sfixed(-0.0582,1,L_SIZE),
				to_sfixed(-0.0578,1,L_SIZE),
				to_sfixed(-0.0574,1,L_SIZE),
				to_sfixed(-0.0571,1,L_SIZE),
				to_sfixed(-0.0567,1,L_SIZE),
				to_sfixed(-0.0563,1,L_SIZE),
				to_sfixed(-0.0560,1,L_SIZE),
				to_sfixed(-0.0556,1,L_SIZE),
				to_sfixed(-0.0552,1,L_SIZE),
				to_sfixed(-0.0549,1,L_SIZE),
				to_sfixed(-0.0545,1,L_SIZE),
				to_sfixed(-0.0541,1,L_SIZE),
				to_sfixed(-0.0538,1,L_SIZE),
				to_sfixed(-0.0534,1,L_SIZE),
				to_sfixed(-0.0531,1,L_SIZE),
				to_sfixed(-0.0527,1,L_SIZE),
				to_sfixed(-0.0523,1,L_SIZE),
				to_sfixed(-0.0520,1,L_SIZE),
				to_sfixed(-0.0516,1,L_SIZE),
				to_sfixed(-0.0512,1,L_SIZE),
				to_sfixed(-0.0509,1,L_SIZE),
				to_sfixed(-0.0505,1,L_SIZE),
				to_sfixed(-0.0501,1,L_SIZE),
				to_sfixed(-0.0498,1,L_SIZE),
				to_sfixed(-0.0494,1,L_SIZE),
				to_sfixed(-0.0490,1,L_SIZE),
				to_sfixed(-0.0487,1,L_SIZE),
				to_sfixed(-0.0483,1,L_SIZE),
				to_sfixed(-0.0479,1,L_SIZE),
				to_sfixed(-0.0476,1,L_SIZE),
				to_sfixed(-0.0472,1,L_SIZE),
				to_sfixed(-0.0468,1,L_SIZE),
				to_sfixed(-0.0465,1,L_SIZE),
				to_sfixed(-0.0461,1,L_SIZE),
				to_sfixed(-0.0457,1,L_SIZE),
				to_sfixed(-0.0454,1,L_SIZE),
				to_sfixed(-0.0450,1,L_SIZE),
				to_sfixed(-0.0446,1,L_SIZE),
				to_sfixed(-0.0443,1,L_SIZE),
				to_sfixed(-0.0439,1,L_SIZE),
				to_sfixed(-0.0436,1,L_SIZE),
				to_sfixed(-0.0432,1,L_SIZE),
				to_sfixed(-0.0428,1,L_SIZE),
				to_sfixed(-0.0425,1,L_SIZE),
				to_sfixed(-0.0421,1,L_SIZE),
				to_sfixed(-0.0417,1,L_SIZE),
				to_sfixed(-0.0414,1,L_SIZE),
				to_sfixed(-0.0410,1,L_SIZE),
				to_sfixed(-0.0406,1,L_SIZE),
				to_sfixed(-0.0403,1,L_SIZE),
				to_sfixed(-0.0399,1,L_SIZE),
				to_sfixed(-0.0395,1,L_SIZE),
				to_sfixed(-0.0392,1,L_SIZE),
				to_sfixed(-0.0388,1,L_SIZE),
				to_sfixed(-0.0384,1,L_SIZE),
				to_sfixed(-0.0381,1,L_SIZE),
				to_sfixed(-0.0377,1,L_SIZE),
				to_sfixed(-0.0373,1,L_SIZE),
				to_sfixed(-0.0370,1,L_SIZE),
				to_sfixed(-0.0366,1,L_SIZE),
				to_sfixed(-0.0362,1,L_SIZE),
				to_sfixed(-0.0359,1,L_SIZE),
				to_sfixed(-0.0355,1,L_SIZE),
				to_sfixed(-0.0351,1,L_SIZE),
				to_sfixed(-0.0348,1,L_SIZE),
				to_sfixed(-0.0344,1,L_SIZE),
				to_sfixed(-0.0340,1,L_SIZE),
				to_sfixed(-0.0337,1,L_SIZE),
				to_sfixed(-0.0333,1,L_SIZE),
				to_sfixed(-0.0329,1,L_SIZE),
				to_sfixed(-0.0326,1,L_SIZE),
				to_sfixed(-0.0322,1,L_SIZE),
				to_sfixed(-0.0318,1,L_SIZE),
				to_sfixed(-0.0315,1,L_SIZE),
				to_sfixed(-0.0311,1,L_SIZE),
				to_sfixed(-0.0308,1,L_SIZE),
				to_sfixed(-0.0304,1,L_SIZE),
				to_sfixed(-0.0300,1,L_SIZE),
				to_sfixed(-0.0297,1,L_SIZE),
				to_sfixed(-0.0293,1,L_SIZE),
				to_sfixed(-0.0289,1,L_SIZE),
				to_sfixed(-0.0286,1,L_SIZE),
				to_sfixed(-0.0282,1,L_SIZE),
				to_sfixed(-0.0278,1,L_SIZE),
				to_sfixed(-0.0275,1,L_SIZE),
				to_sfixed(-0.0271,1,L_SIZE),
				to_sfixed(-0.0267,1,L_SIZE),
				to_sfixed(-0.0264,1,L_SIZE),
				to_sfixed(-0.0260,1,L_SIZE),
				to_sfixed(-0.0256,1,L_SIZE),
				to_sfixed(-0.0253,1,L_SIZE),
				to_sfixed(-0.0249,1,L_SIZE),
				to_sfixed(-0.0245,1,L_SIZE),
				to_sfixed(-0.0242,1,L_SIZE),
				to_sfixed(-0.0238,1,L_SIZE),
				to_sfixed(-0.0234,1,L_SIZE),
				to_sfixed(-0.0231,1,L_SIZE),
				to_sfixed(-0.0227,1,L_SIZE),
				to_sfixed(-0.0223,1,L_SIZE),
				to_sfixed(-0.0220,1,L_SIZE),
				to_sfixed(-0.0216,1,L_SIZE),
				to_sfixed(-0.0212,1,L_SIZE),
				to_sfixed(-0.0209,1,L_SIZE),
				to_sfixed(-0.0205,1,L_SIZE),
				to_sfixed(-0.0201,1,L_SIZE),
				to_sfixed(-0.0198,1,L_SIZE),
				to_sfixed(-0.0194,1,L_SIZE),
				to_sfixed(-0.0190,1,L_SIZE),
				to_sfixed(-0.0187,1,L_SIZE),
				to_sfixed(-0.0183,1,L_SIZE),
				to_sfixed(-0.0179,1,L_SIZE),
				to_sfixed(-0.0176,1,L_SIZE),
				to_sfixed(-0.0172,1,L_SIZE),
				to_sfixed(-0.0168,1,L_SIZE),
				to_sfixed(-0.0165,1,L_SIZE),
				to_sfixed(-0.0161,1,L_SIZE),
				to_sfixed(-0.0157,1,L_SIZE),
				to_sfixed(-0.0154,1,L_SIZE),
				to_sfixed(-0.0150,1,L_SIZE),
				to_sfixed(-0.0146,1,L_SIZE),
				to_sfixed(-0.0143,1,L_SIZE),
				to_sfixed(-0.0139,1,L_SIZE),
				to_sfixed(-0.0135,1,L_SIZE),
				to_sfixed(-0.0132,1,L_SIZE),
				to_sfixed(-0.0128,1,L_SIZE),
				to_sfixed(-0.0125,1,L_SIZE),
				to_sfixed(-0.0121,1,L_SIZE),
				to_sfixed(-0.0117,1,L_SIZE),
				to_sfixed(-0.0114,1,L_SIZE),
				to_sfixed(-0.0110,1,L_SIZE),
				to_sfixed(-0.0106,1,L_SIZE),
				to_sfixed(-0.0103,1,L_SIZE),
				to_sfixed(-0.0099,1,L_SIZE),
				to_sfixed(-0.0095,1,L_SIZE),
				to_sfixed(-0.0092,1,L_SIZE),
				to_sfixed(-0.0088,1,L_SIZE),
				to_sfixed(-0.0084,1,L_SIZE),
				to_sfixed(-0.0081,1,L_SIZE),
				to_sfixed(-0.0077,1,L_SIZE),
				to_sfixed(-0.0073,1,L_SIZE),
				to_sfixed(-0.0070,1,L_SIZE),
				to_sfixed(-0.0066,1,L_SIZE),
				to_sfixed(-0.0062,1,L_SIZE),
				to_sfixed(-0.0059,1,L_SIZE),
				to_sfixed(-0.0055,1,L_SIZE),
				to_sfixed(-0.0051,1,L_SIZE),
				to_sfixed(-0.0048,1,L_SIZE),
				to_sfixed(-0.0044,1,L_SIZE),
				to_sfixed(-0.0040,1,L_SIZE),
				to_sfixed(-0.0037,1,L_SIZE),
				to_sfixed(-0.0033,1,L_SIZE),
				to_sfixed(-0.0029,1,L_SIZE),
				to_sfixed(-0.0026,1,L_SIZE),
				to_sfixed(-0.0022,1,L_SIZE),
				to_sfixed(-0.0018,1,L_SIZE),
				to_sfixed(-0.0015,1,L_SIZE),
				to_sfixed(-0.0011,1,L_SIZE),
				to_sfixed(-0.0007,1,L_SIZE),
				to_sfixed(-0.0004,1,L_SIZE),
				to_sfixed(0.0000,1,L_SIZE),
				to_sfixed(0.0004,1,L_SIZE),
				to_sfixed(0.0007,1,L_SIZE),
				to_sfixed(0.0011,1,L_SIZE),
				to_sfixed(0.0015,1,L_SIZE),
				to_sfixed(0.0018,1,L_SIZE),
				to_sfixed(0.0022,1,L_SIZE),
				to_sfixed(0.0026,1,L_SIZE),
				to_sfixed(0.0029,1,L_SIZE),
				to_sfixed(0.0033,1,L_SIZE),
				to_sfixed(0.0037,1,L_SIZE),
				to_sfixed(0.0040,1,L_SIZE),
				to_sfixed(0.0044,1,L_SIZE),
				to_sfixed(0.0048,1,L_SIZE),
				to_sfixed(0.0051,1,L_SIZE),
				to_sfixed(0.0055,1,L_SIZE),
				to_sfixed(0.0059,1,L_SIZE),
				to_sfixed(0.0062,1,L_SIZE),
				to_sfixed(0.0066,1,L_SIZE),
				to_sfixed(0.0070,1,L_SIZE),
				to_sfixed(0.0073,1,L_SIZE),
				to_sfixed(0.0077,1,L_SIZE),
				to_sfixed(0.0081,1,L_SIZE),
				to_sfixed(0.0084,1,L_SIZE),
				to_sfixed(0.0088,1,L_SIZE),
				to_sfixed(0.0092,1,L_SIZE),
				to_sfixed(0.0095,1,L_SIZE),
				to_sfixed(0.0099,1,L_SIZE),
				to_sfixed(0.0103,1,L_SIZE),
				to_sfixed(0.0106,1,L_SIZE),
				to_sfixed(0.0110,1,L_SIZE),
				to_sfixed(0.0114,1,L_SIZE),
				to_sfixed(0.0117,1,L_SIZE),
				to_sfixed(0.0121,1,L_SIZE),
				to_sfixed(0.0125,1,L_SIZE),
				to_sfixed(0.0128,1,L_SIZE),
				to_sfixed(0.0132,1,L_SIZE),
				to_sfixed(0.0135,1,L_SIZE),
				to_sfixed(0.0139,1,L_SIZE),
				to_sfixed(0.0143,1,L_SIZE),
				to_sfixed(0.0146,1,L_SIZE),
				to_sfixed(0.0150,1,L_SIZE),
				to_sfixed(0.0154,1,L_SIZE),
				to_sfixed(0.0157,1,L_SIZE),
				to_sfixed(0.0161,1,L_SIZE),
				to_sfixed(0.0165,1,L_SIZE),
				to_sfixed(0.0168,1,L_SIZE),
				to_sfixed(0.0172,1,L_SIZE),
				to_sfixed(0.0176,1,L_SIZE),
				to_sfixed(0.0179,1,L_SIZE),
				to_sfixed(0.0183,1,L_SIZE),
				to_sfixed(0.0187,1,L_SIZE),
				to_sfixed(0.0190,1,L_SIZE),
				to_sfixed(0.0194,1,L_SIZE),
				to_sfixed(0.0198,1,L_SIZE),
				to_sfixed(0.0201,1,L_SIZE),
				to_sfixed(0.0205,1,L_SIZE),
				to_sfixed(0.0209,1,L_SIZE),
				to_sfixed(0.0212,1,L_SIZE),
				to_sfixed(0.0216,1,L_SIZE),
				to_sfixed(0.0220,1,L_SIZE),
				to_sfixed(0.0223,1,L_SIZE),
				to_sfixed(0.0227,1,L_SIZE),
				to_sfixed(0.0231,1,L_SIZE),
				to_sfixed(0.0234,1,L_SIZE),
				to_sfixed(0.0238,1,L_SIZE),
				to_sfixed(0.0242,1,L_SIZE),
				to_sfixed(0.0245,1,L_SIZE),
				to_sfixed(0.0249,1,L_SIZE),
				to_sfixed(0.0253,1,L_SIZE),
				to_sfixed(0.0256,1,L_SIZE),
				to_sfixed(0.0260,1,L_SIZE),
				to_sfixed(0.0264,1,L_SIZE),
				to_sfixed(0.0267,1,L_SIZE),
				to_sfixed(0.0271,1,L_SIZE),
				to_sfixed(0.0275,1,L_SIZE),
				to_sfixed(0.0278,1,L_SIZE),
				to_sfixed(0.0282,1,L_SIZE),
				to_sfixed(0.0286,1,L_SIZE),
				to_sfixed(0.0289,1,L_SIZE),
				to_sfixed(0.0293,1,L_SIZE),
				to_sfixed(0.0297,1,L_SIZE),
				to_sfixed(0.0300,1,L_SIZE),
				to_sfixed(0.0304,1,L_SIZE),
				to_sfixed(0.0308,1,L_SIZE),
				to_sfixed(0.0311,1,L_SIZE),
				to_sfixed(0.0315,1,L_SIZE),
				to_sfixed(0.0318,1,L_SIZE),
				to_sfixed(0.0322,1,L_SIZE),
				to_sfixed(0.0326,1,L_SIZE),
				to_sfixed(0.0329,1,L_SIZE),
				to_sfixed(0.0333,1,L_SIZE),
				to_sfixed(0.0337,1,L_SIZE),
				to_sfixed(0.0340,1,L_SIZE),
				to_sfixed(0.0344,1,L_SIZE),
				to_sfixed(0.0348,1,L_SIZE),
				to_sfixed(0.0351,1,L_SIZE),
				to_sfixed(0.0355,1,L_SIZE),
				to_sfixed(0.0359,1,L_SIZE),
				to_sfixed(0.0362,1,L_SIZE),
				to_sfixed(0.0366,1,L_SIZE),
				to_sfixed(0.0370,1,L_SIZE),
				to_sfixed(0.0373,1,L_SIZE),
				to_sfixed(0.0377,1,L_SIZE),
				to_sfixed(0.0381,1,L_SIZE),
				to_sfixed(0.0384,1,L_SIZE),
				to_sfixed(0.0388,1,L_SIZE),
				to_sfixed(0.0392,1,L_SIZE),
				to_sfixed(0.0395,1,L_SIZE),
				to_sfixed(0.0399,1,L_SIZE),
				to_sfixed(0.0403,1,L_SIZE),
				to_sfixed(0.0406,1,L_SIZE),
				to_sfixed(0.0410,1,L_SIZE),
				to_sfixed(0.0414,1,L_SIZE),
				to_sfixed(0.0417,1,L_SIZE),
				to_sfixed(0.0421,1,L_SIZE),
				to_sfixed(0.0425,1,L_SIZE),
				to_sfixed(0.0428,1,L_SIZE),
				to_sfixed(0.0432,1,L_SIZE),
				to_sfixed(0.0436,1,L_SIZE),
				to_sfixed(0.0439,1,L_SIZE),
				to_sfixed(0.0443,1,L_SIZE),
				to_sfixed(0.0446,1,L_SIZE),
				to_sfixed(0.0450,1,L_SIZE),
				to_sfixed(0.0454,1,L_SIZE),
				to_sfixed(0.0457,1,L_SIZE),
				to_sfixed(0.0461,1,L_SIZE),
				to_sfixed(0.0465,1,L_SIZE),
				to_sfixed(0.0468,1,L_SIZE),
				to_sfixed(0.0472,1,L_SIZE),
				to_sfixed(0.0476,1,L_SIZE),
				to_sfixed(0.0479,1,L_SIZE),
				to_sfixed(0.0483,1,L_SIZE),
				to_sfixed(0.0487,1,L_SIZE),
				to_sfixed(0.0490,1,L_SIZE),
				to_sfixed(0.0494,1,L_SIZE),
				to_sfixed(0.0498,1,L_SIZE),
				to_sfixed(0.0501,1,L_SIZE),
				to_sfixed(0.0505,1,L_SIZE),
				to_sfixed(0.0509,1,L_SIZE),
				to_sfixed(0.0512,1,L_SIZE),
				to_sfixed(0.0516,1,L_SIZE),
				to_sfixed(0.0520,1,L_SIZE),
				to_sfixed(0.0523,1,L_SIZE),
				to_sfixed(0.0527,1,L_SIZE),
				to_sfixed(0.0531,1,L_SIZE),
				to_sfixed(0.0534,1,L_SIZE),
				to_sfixed(0.0538,1,L_SIZE),
				to_sfixed(0.0541,1,L_SIZE),
				to_sfixed(0.0545,1,L_SIZE),
				to_sfixed(0.0549,1,L_SIZE),
				to_sfixed(0.0552,1,L_SIZE),
				to_sfixed(0.0556,1,L_SIZE),
				to_sfixed(0.0560,1,L_SIZE),
				to_sfixed(0.0563,1,L_SIZE),
				to_sfixed(0.0567,1,L_SIZE),
				to_sfixed(0.0571,1,L_SIZE),
				to_sfixed(0.0574,1,L_SIZE),
				to_sfixed(0.0578,1,L_SIZE),
				to_sfixed(0.0582,1,L_SIZE),
				to_sfixed(0.0585,1,L_SIZE),
				to_sfixed(0.0589,1,L_SIZE),
				to_sfixed(0.0593,1,L_SIZE),
				to_sfixed(0.0596,1,L_SIZE),
				to_sfixed(0.0600,1,L_SIZE),
				to_sfixed(0.0604,1,L_SIZE),
				to_sfixed(0.0607,1,L_SIZE),
				to_sfixed(0.0611,1,L_SIZE),
				to_sfixed(0.0614,1,L_SIZE),
				to_sfixed(0.0618,1,L_SIZE),
				to_sfixed(0.0622,1,L_SIZE),
				to_sfixed(0.0625,1,L_SIZE),
				to_sfixed(0.0629,1,L_SIZE),
				to_sfixed(0.0633,1,L_SIZE),
				to_sfixed(0.0636,1,L_SIZE),
				to_sfixed(0.0640,1,L_SIZE),
				to_sfixed(0.0644,1,L_SIZE),
				to_sfixed(0.0647,1,L_SIZE),
				to_sfixed(0.0651,1,L_SIZE),
				to_sfixed(0.0655,1,L_SIZE),
				to_sfixed(0.0658,1,L_SIZE),
				to_sfixed(0.0662,1,L_SIZE),
				to_sfixed(0.0666,1,L_SIZE),
				to_sfixed(0.0669,1,L_SIZE),
				to_sfixed(0.0673,1,L_SIZE),
				to_sfixed(0.0676,1,L_SIZE),
				to_sfixed(0.0680,1,L_SIZE),
				to_sfixed(0.0684,1,L_SIZE),
				to_sfixed(0.0687,1,L_SIZE),
				to_sfixed(0.0691,1,L_SIZE),
				to_sfixed(0.0695,1,L_SIZE),
				to_sfixed(0.0698,1,L_SIZE),
				to_sfixed(0.0702,1,L_SIZE),
				to_sfixed(0.0706,1,L_SIZE),
				to_sfixed(0.0709,1,L_SIZE),
				to_sfixed(0.0713,1,L_SIZE),
				to_sfixed(0.0717,1,L_SIZE),
				to_sfixed(0.0720,1,L_SIZE),
				to_sfixed(0.0724,1,L_SIZE),
				to_sfixed(0.0727,1,L_SIZE),
				to_sfixed(0.0731,1,L_SIZE),
				to_sfixed(0.0735,1,L_SIZE),
				to_sfixed(0.0738,1,L_SIZE),
				to_sfixed(0.0742,1,L_SIZE),
				to_sfixed(0.0746,1,L_SIZE),
				to_sfixed(0.0749,1,L_SIZE),
				to_sfixed(0.0753,1,L_SIZE),
				to_sfixed(0.0757,1,L_SIZE),
				to_sfixed(0.0760,1,L_SIZE),
				to_sfixed(0.0764,1,L_SIZE),
				to_sfixed(0.0768,1,L_SIZE),
				to_sfixed(0.0771,1,L_SIZE),
				to_sfixed(0.0775,1,L_SIZE),
				to_sfixed(0.0778,1,L_SIZE),
				to_sfixed(0.0782,1,L_SIZE),
				to_sfixed(0.0786,1,L_SIZE),
				to_sfixed(0.0789,1,L_SIZE),
				to_sfixed(0.0793,1,L_SIZE),
				to_sfixed(0.0797,1,L_SIZE),
				to_sfixed(0.0800,1,L_SIZE),
				to_sfixed(0.0804,1,L_SIZE),
				to_sfixed(0.0808,1,L_SIZE),
				to_sfixed(0.0811,1,L_SIZE),
				to_sfixed(0.0815,1,L_SIZE),
				to_sfixed(0.0818,1,L_SIZE),
				to_sfixed(0.0822,1,L_SIZE),
				to_sfixed(0.0826,1,L_SIZE),
				to_sfixed(0.0829,1,L_SIZE),
				to_sfixed(0.0833,1,L_SIZE),
				to_sfixed(0.0837,1,L_SIZE),
				to_sfixed(0.0840,1,L_SIZE),
				to_sfixed(0.0844,1,L_SIZE),
				to_sfixed(0.0848,1,L_SIZE),
				to_sfixed(0.0851,1,L_SIZE),
				to_sfixed(0.0855,1,L_SIZE),
				to_sfixed(0.0858,1,L_SIZE),
				to_sfixed(0.0862,1,L_SIZE),
				to_sfixed(0.0866,1,L_SIZE),
				to_sfixed(0.0869,1,L_SIZE),
				to_sfixed(0.0873,1,L_SIZE),
				to_sfixed(0.0877,1,L_SIZE),
				to_sfixed(0.0880,1,L_SIZE),
				to_sfixed(0.0884,1,L_SIZE),
				to_sfixed(0.0888,1,L_SIZE),
				to_sfixed(0.0891,1,L_SIZE),
				to_sfixed(0.0895,1,L_SIZE),
				to_sfixed(0.0898,1,L_SIZE),
				to_sfixed(0.0902,1,L_SIZE),
				to_sfixed(0.0906,1,L_SIZE),
				to_sfixed(0.0909,1,L_SIZE),
				to_sfixed(0.0913,1,L_SIZE),
				to_sfixed(0.0917,1,L_SIZE),
				to_sfixed(0.0920,1,L_SIZE),
				to_sfixed(0.0924,1,L_SIZE),
				to_sfixed(0.0928,1,L_SIZE),
				to_sfixed(0.0931,1,L_SIZE),
				to_sfixed(0.0935,1,L_SIZE),
				to_sfixed(0.0938,1,L_SIZE),
				to_sfixed(0.0942,1,L_SIZE),
				to_sfixed(0.0946,1,L_SIZE),
				to_sfixed(0.0949,1,L_SIZE),
				to_sfixed(0.0953,1,L_SIZE),
				to_sfixed(0.0957,1,L_SIZE),
				to_sfixed(0.0960,1,L_SIZE),
				to_sfixed(0.0964,1,L_SIZE),
				to_sfixed(0.0967,1,L_SIZE),
				to_sfixed(0.0971,1,L_SIZE),
				to_sfixed(0.0975,1,L_SIZE),
				to_sfixed(0.0978,1,L_SIZE),
				to_sfixed(0.0982,1,L_SIZE),
				to_sfixed(0.0986,1,L_SIZE),
				to_sfixed(0.0989,1,L_SIZE),
				to_sfixed(0.0993,1,L_SIZE),
				to_sfixed(0.0996,1,L_SIZE),
				to_sfixed(0.1000,1,L_SIZE),
				to_sfixed(0.1004,1,L_SIZE),
				to_sfixed(0.1007,1,L_SIZE),
				to_sfixed(0.1011,1,L_SIZE),
				to_sfixed(0.1015,1,L_SIZE),
				to_sfixed(0.1018,1,L_SIZE),
				to_sfixed(0.1022,1,L_SIZE),
				to_sfixed(0.1025,1,L_SIZE),
				to_sfixed(0.1029,1,L_SIZE),
				to_sfixed(0.1033,1,L_SIZE),
				to_sfixed(0.1036,1,L_SIZE),
				to_sfixed(0.1040,1,L_SIZE),
				to_sfixed(0.1044,1,L_SIZE),
				to_sfixed(0.1047,1,L_SIZE),
				to_sfixed(0.1051,1,L_SIZE),
				to_sfixed(0.1054,1,L_SIZE),
				to_sfixed(0.1058,1,L_SIZE),
				to_sfixed(0.1062,1,L_SIZE),
				to_sfixed(0.1065,1,L_SIZE),
				to_sfixed(0.1069,1,L_SIZE),
				to_sfixed(0.1073,1,L_SIZE),
				to_sfixed(0.1076,1,L_SIZE),
				to_sfixed(0.1080,1,L_SIZE),
				to_sfixed(0.1083,1,L_SIZE),
				to_sfixed(0.1087,1,L_SIZE),
				to_sfixed(0.1091,1,L_SIZE),
				to_sfixed(0.1094,1,L_SIZE),
				to_sfixed(0.1098,1,L_SIZE),
				to_sfixed(0.1101,1,L_SIZE),
				to_sfixed(0.1105,1,L_SIZE),
				to_sfixed(0.1109,1,L_SIZE),
				to_sfixed(0.1112,1,L_SIZE),
				to_sfixed(0.1116,1,L_SIZE),
				to_sfixed(0.1120,1,L_SIZE),
				to_sfixed(0.1123,1,L_SIZE),
				to_sfixed(0.1127,1,L_SIZE),
				to_sfixed(0.1130,1,L_SIZE),
				to_sfixed(0.1134,1,L_SIZE),
				to_sfixed(0.1138,1,L_SIZE),
				to_sfixed(0.1141,1,L_SIZE),
				to_sfixed(0.1145,1,L_SIZE),
				to_sfixed(0.1148,1,L_SIZE),
				to_sfixed(0.1152,1,L_SIZE),
				to_sfixed(0.1156,1,L_SIZE),
				to_sfixed(0.1159,1,L_SIZE),
				to_sfixed(0.1163,1,L_SIZE),
				to_sfixed(0.1167,1,L_SIZE),
				to_sfixed(0.1170,1,L_SIZE),
				to_sfixed(0.1174,1,L_SIZE),
				to_sfixed(0.1177,1,L_SIZE),
				to_sfixed(0.1181,1,L_SIZE),
				to_sfixed(0.1185,1,L_SIZE),
				to_sfixed(0.1188,1,L_SIZE),
				to_sfixed(0.1192,1,L_SIZE),
				to_sfixed(0.1195,1,L_SIZE),
				to_sfixed(0.1199,1,L_SIZE),
				to_sfixed(0.1203,1,L_SIZE),
				to_sfixed(0.1206,1,L_SIZE),
				to_sfixed(0.1210,1,L_SIZE),
				to_sfixed(0.1213,1,L_SIZE),
				to_sfixed(0.1217,1,L_SIZE),
				to_sfixed(0.1221,1,L_SIZE),
				to_sfixed(0.1224,1,L_SIZE),
				to_sfixed(0.1228,1,L_SIZE),
				to_sfixed(0.1232,1,L_SIZE),
				to_sfixed(0.1235,1,L_SIZE),
				to_sfixed(0.1239,1,L_SIZE),
				to_sfixed(0.1242,1,L_SIZE),
				to_sfixed(0.1246,1,L_SIZE),
				to_sfixed(0.1250,1,L_SIZE),
				to_sfixed(0.1253,1,L_SIZE),
				to_sfixed(0.1257,1,L_SIZE),
				to_sfixed(0.1260,1,L_SIZE),
				to_sfixed(0.1264,1,L_SIZE),
				to_sfixed(0.1268,1,L_SIZE),
				to_sfixed(0.1271,1,L_SIZE),
				to_sfixed(0.1275,1,L_SIZE),
				to_sfixed(0.1278,1,L_SIZE),
				to_sfixed(0.1282,1,L_SIZE),
				to_sfixed(0.1286,1,L_SIZE),
				to_sfixed(0.1289,1,L_SIZE),
				to_sfixed(0.1293,1,L_SIZE),
				to_sfixed(0.1296,1,L_SIZE),
				to_sfixed(0.1300,1,L_SIZE),
				to_sfixed(0.1304,1,L_SIZE),
				to_sfixed(0.1307,1,L_SIZE),
				to_sfixed(0.1311,1,L_SIZE),
				to_sfixed(0.1314,1,L_SIZE),
				to_sfixed(0.1318,1,L_SIZE),
				to_sfixed(0.1322,1,L_SIZE),
				to_sfixed(0.1325,1,L_SIZE),
				to_sfixed(0.1329,1,L_SIZE),
				to_sfixed(0.1332,1,L_SIZE),
				to_sfixed(0.1336,1,L_SIZE),
				to_sfixed(0.1340,1,L_SIZE),
				to_sfixed(0.1343,1,L_SIZE),
				to_sfixed(0.1347,1,L_SIZE),
				to_sfixed(0.1350,1,L_SIZE),
				to_sfixed(0.1354,1,L_SIZE),
				to_sfixed(0.1358,1,L_SIZE),
				to_sfixed(0.1361,1,L_SIZE),
				to_sfixed(0.1365,1,L_SIZE),
				to_sfixed(0.1368,1,L_SIZE),
				to_sfixed(0.1372,1,L_SIZE),
				to_sfixed(0.1376,1,L_SIZE),
				to_sfixed(0.1379,1,L_SIZE),
				to_sfixed(0.1383,1,L_SIZE),
				to_sfixed(0.1386,1,L_SIZE),
				to_sfixed(0.1390,1,L_SIZE),
				to_sfixed(0.1393,1,L_SIZE),
				to_sfixed(0.1397,1,L_SIZE),
				to_sfixed(0.1401,1,L_SIZE),
				to_sfixed(0.1404,1,L_SIZE),
				to_sfixed(0.1408,1,L_SIZE),
				to_sfixed(0.1411,1,L_SIZE),
				to_sfixed(0.1415,1,L_SIZE),
				to_sfixed(0.1419,1,L_SIZE),
				to_sfixed(0.1422,1,L_SIZE),
				to_sfixed(0.1426,1,L_SIZE),
				to_sfixed(0.1429,1,L_SIZE),
				to_sfixed(0.1433,1,L_SIZE),
				to_sfixed(0.1437,1,L_SIZE),
				to_sfixed(0.1440,1,L_SIZE),
				to_sfixed(0.1444,1,L_SIZE),
				to_sfixed(0.1447,1,L_SIZE),
				to_sfixed(0.1451,1,L_SIZE),
				to_sfixed(0.1454,1,L_SIZE),
				to_sfixed(0.1458,1,L_SIZE),
				to_sfixed(0.1462,1,L_SIZE),
				to_sfixed(0.1465,1,L_SIZE),
				to_sfixed(0.1469,1,L_SIZE),
				to_sfixed(0.1472,1,L_SIZE),
				to_sfixed(0.1476,1,L_SIZE),
				to_sfixed(0.1480,1,L_SIZE),
				to_sfixed(0.1483,1,L_SIZE),
				to_sfixed(0.1487,1,L_SIZE),
				to_sfixed(0.1490,1,L_SIZE),
				to_sfixed(0.1494,1,L_SIZE),
				to_sfixed(0.1497,1,L_SIZE),
				to_sfixed(0.1501,1,L_SIZE),
				to_sfixed(0.1505,1,L_SIZE),
				to_sfixed(0.1508,1,L_SIZE),
				to_sfixed(0.1512,1,L_SIZE),
				to_sfixed(0.1515,1,L_SIZE),
				to_sfixed(0.1519,1,L_SIZE),
				to_sfixed(0.1522,1,L_SIZE),
				to_sfixed(0.1526,1,L_SIZE),
				to_sfixed(0.1530,1,L_SIZE),
				to_sfixed(0.1533,1,L_SIZE),
				to_sfixed(0.1537,1,L_SIZE),
				to_sfixed(0.1540,1,L_SIZE),
				to_sfixed(0.1544,1,L_SIZE),
				to_sfixed(0.1548,1,L_SIZE),
				to_sfixed(0.1551,1,L_SIZE),
				to_sfixed(0.1555,1,L_SIZE),
				to_sfixed(0.1558,1,L_SIZE),
				to_sfixed(0.1562,1,L_SIZE),
				to_sfixed(0.1565,1,L_SIZE),
				to_sfixed(0.1569,1,L_SIZE),
				to_sfixed(0.1573,1,L_SIZE),
				to_sfixed(0.1576,1,L_SIZE),
				to_sfixed(0.1580,1,L_SIZE),
				to_sfixed(0.1583,1,L_SIZE),
				to_sfixed(0.1587,1,L_SIZE),
				to_sfixed(0.1590,1,L_SIZE),
				to_sfixed(0.1594,1,L_SIZE),
				to_sfixed(0.1598,1,L_SIZE),
				to_sfixed(0.1601,1,L_SIZE),
				to_sfixed(0.1605,1,L_SIZE),
				to_sfixed(0.1608,1,L_SIZE),
				to_sfixed(0.1612,1,L_SIZE),
				to_sfixed(0.1615,1,L_SIZE),
				to_sfixed(0.1619,1,L_SIZE),
				to_sfixed(0.1622,1,L_SIZE),
				to_sfixed(0.1626,1,L_SIZE),
				to_sfixed(0.1630,1,L_SIZE),
				to_sfixed(0.1633,1,L_SIZE),
				to_sfixed(0.1637,1,L_SIZE),
				to_sfixed(0.1640,1,L_SIZE),
				to_sfixed(0.1644,1,L_SIZE),
				to_sfixed(0.1647,1,L_SIZE),
				to_sfixed(0.1651,1,L_SIZE),
				to_sfixed(0.1655,1,L_SIZE),
				to_sfixed(0.1658,1,L_SIZE),
				to_sfixed(0.1662,1,L_SIZE),
				to_sfixed(0.1665,1,L_SIZE),
				to_sfixed(0.1669,1,L_SIZE),
				to_sfixed(0.1672,1,L_SIZE),
				to_sfixed(0.1676,1,L_SIZE),
				to_sfixed(0.1679,1,L_SIZE),
				to_sfixed(0.1683,1,L_SIZE),
				to_sfixed(0.1687,1,L_SIZE),
				to_sfixed(0.1690,1,L_SIZE),
				to_sfixed(0.1694,1,L_SIZE),
				to_sfixed(0.1697,1,L_SIZE),
				to_sfixed(0.1701,1,L_SIZE),
				to_sfixed(0.1704,1,L_SIZE),
				to_sfixed(0.1708,1,L_SIZE),
				to_sfixed(0.1712,1,L_SIZE),
				to_sfixed(0.1715,1,L_SIZE),
				to_sfixed(0.1719,1,L_SIZE),
				to_sfixed(0.1722,1,L_SIZE),
				to_sfixed(0.1726,1,L_SIZE),
				to_sfixed(0.1729,1,L_SIZE),
				to_sfixed(0.1733,1,L_SIZE),
				to_sfixed(0.1736,1,L_SIZE),
				to_sfixed(0.1740,1,L_SIZE),
				to_sfixed(0.1743,1,L_SIZE),
				to_sfixed(0.1747,1,L_SIZE),
				to_sfixed(0.1751,1,L_SIZE),
				to_sfixed(0.1754,1,L_SIZE),
				to_sfixed(0.1758,1,L_SIZE),
				to_sfixed(0.1761,1,L_SIZE),
				to_sfixed(0.1765,1,L_SIZE),
				to_sfixed(0.1768,1,L_SIZE),
				to_sfixed(0.1772,1,L_SIZE),
				to_sfixed(0.1775,1,L_SIZE),
				to_sfixed(0.1779,1,L_SIZE),
				to_sfixed(0.1783,1,L_SIZE),
				to_sfixed(0.1786,1,L_SIZE),
				to_sfixed(0.1790,1,L_SIZE),
				to_sfixed(0.1793,1,L_SIZE),
				to_sfixed(0.1797,1,L_SIZE),
				to_sfixed(0.1800,1,L_SIZE),
				to_sfixed(0.1804,1,L_SIZE),
				to_sfixed(0.1807,1,L_SIZE),
				to_sfixed(0.1811,1,L_SIZE),
				to_sfixed(0.1814,1,L_SIZE),
				to_sfixed(0.1818,1,L_SIZE),
				to_sfixed(0.1821,1,L_SIZE),
				to_sfixed(0.1825,1,L_SIZE),
				to_sfixed(0.1829,1,L_SIZE),
				to_sfixed(0.1832,1,L_SIZE),
				to_sfixed(0.1836,1,L_SIZE),
				to_sfixed(0.1839,1,L_SIZE),
				to_sfixed(0.1843,1,L_SIZE),
				to_sfixed(0.1846,1,L_SIZE),
				to_sfixed(0.1850,1,L_SIZE),
				to_sfixed(0.1853,1,L_SIZE),
				to_sfixed(0.1857,1,L_SIZE),
				to_sfixed(0.1860,1,L_SIZE),
				to_sfixed(0.1864,1,L_SIZE),
				to_sfixed(0.1867,1,L_SIZE),
				to_sfixed(0.1871,1,L_SIZE),
				to_sfixed(0.1875,1,L_SIZE),
				to_sfixed(0.1878,1,L_SIZE),
				to_sfixed(0.1882,1,L_SIZE),
				to_sfixed(0.1885,1,L_SIZE),
				to_sfixed(0.1889,1,L_SIZE),
				to_sfixed(0.1892,1,L_SIZE),
				to_sfixed(0.1896,1,L_SIZE),
				to_sfixed(0.1899,1,L_SIZE),
				to_sfixed(0.1903,1,L_SIZE),
				to_sfixed(0.1906,1,L_SIZE),
				to_sfixed(0.1910,1,L_SIZE),
				to_sfixed(0.1913,1,L_SIZE),
				to_sfixed(0.1917,1,L_SIZE),
				to_sfixed(0.1920,1,L_SIZE),
				to_sfixed(0.1924,1,L_SIZE),
				to_sfixed(0.1927,1,L_SIZE),
				to_sfixed(0.1931,1,L_SIZE),
				to_sfixed(0.1935,1,L_SIZE),
				to_sfixed(0.1938,1,L_SIZE),
				to_sfixed(0.1942,1,L_SIZE),
				to_sfixed(0.1945,1,L_SIZE),
				to_sfixed(0.1949,1,L_SIZE),
				to_sfixed(0.1952,1,L_SIZE),
				to_sfixed(0.1956,1,L_SIZE),
				to_sfixed(0.1959,1,L_SIZE),
				to_sfixed(0.1963,1,L_SIZE),
				to_sfixed(0.1966,1,L_SIZE),
				to_sfixed(0.1970,1,L_SIZE),
				to_sfixed(0.1973,1,L_SIZE),
				to_sfixed(0.1977,1,L_SIZE),
				to_sfixed(0.1980,1,L_SIZE),
				to_sfixed(0.1984,1,L_SIZE),
				to_sfixed(0.1987,1,L_SIZE),
				to_sfixed(0.1991,1,L_SIZE),
				to_sfixed(0.1994,1,L_SIZE),
				to_sfixed(0.1998,1,L_SIZE),
				to_sfixed(0.2001,1,L_SIZE),
				to_sfixed(0.2005,1,L_SIZE),
				to_sfixed(0.2008,1,L_SIZE),
				to_sfixed(0.2012,1,L_SIZE),
				to_sfixed(0.2015,1,L_SIZE),
				to_sfixed(0.2019,1,L_SIZE),
				to_sfixed(0.2023,1,L_SIZE),
				to_sfixed(0.2026,1,L_SIZE),
				to_sfixed(0.2030,1,L_SIZE),
				to_sfixed(0.2033,1,L_SIZE),
				to_sfixed(0.2037,1,L_SIZE),
				to_sfixed(0.2040,1,L_SIZE),
				to_sfixed(0.2044,1,L_SIZE),
				to_sfixed(0.2047,1,L_SIZE),
				to_sfixed(0.2051,1,L_SIZE),
				to_sfixed(0.2054,1,L_SIZE),
				to_sfixed(0.2058,1,L_SIZE),
				to_sfixed(0.2061,1,L_SIZE),
				to_sfixed(0.2065,1,L_SIZE),
				to_sfixed(0.2068,1,L_SIZE),
				to_sfixed(0.2072,1,L_SIZE),
				to_sfixed(0.2075,1,L_SIZE),
				to_sfixed(0.2079,1,L_SIZE),
				to_sfixed(0.2082,1,L_SIZE),
				to_sfixed(0.2086,1,L_SIZE),
				to_sfixed(0.2089,1,L_SIZE),
				to_sfixed(0.2093,1,L_SIZE),
				to_sfixed(0.2096,1,L_SIZE),
				to_sfixed(0.2100,1,L_SIZE),
				to_sfixed(0.2103,1,L_SIZE),
				to_sfixed(0.2107,1,L_SIZE),
				to_sfixed(0.2110,1,L_SIZE),
				to_sfixed(0.2114,1,L_SIZE),
				to_sfixed(0.2117,1,L_SIZE),
				to_sfixed(0.2121,1,L_SIZE),
				to_sfixed(0.2124,1,L_SIZE),
				to_sfixed(0.2128,1,L_SIZE),
				to_sfixed(0.2131,1,L_SIZE),
				to_sfixed(0.2135,1,L_SIZE),
				to_sfixed(0.2138,1,L_SIZE),
				to_sfixed(0.2142,1,L_SIZE),
				to_sfixed(0.2145,1,L_SIZE),
				to_sfixed(0.2149,1,L_SIZE),
				to_sfixed(0.2152,1,L_SIZE),
				to_sfixed(0.2156,1,L_SIZE),
				to_sfixed(0.2159,1,L_SIZE),
				to_sfixed(0.2163,1,L_SIZE),
				to_sfixed(0.2166,1,L_SIZE),
				to_sfixed(0.2170,1,L_SIZE),
				to_sfixed(0.2173,1,L_SIZE),
				to_sfixed(0.2177,1,L_SIZE),
				to_sfixed(0.2180,1,L_SIZE),
				to_sfixed(0.2184,1,L_SIZE),
				to_sfixed(0.2187,1,L_SIZE),
				to_sfixed(0.2190,1,L_SIZE),
				to_sfixed(0.2194,1,L_SIZE),
				to_sfixed(0.2197,1,L_SIZE),
				to_sfixed(0.2201,1,L_SIZE),
				to_sfixed(0.2204,1,L_SIZE),
				to_sfixed(0.2208,1,L_SIZE),
				to_sfixed(0.2211,1,L_SIZE),
				to_sfixed(0.2215,1,L_SIZE),
				to_sfixed(0.2218,1,L_SIZE),
				to_sfixed(0.2222,1,L_SIZE),
				to_sfixed(0.2225,1,L_SIZE),
				to_sfixed(0.2229,1,L_SIZE),
				to_sfixed(0.2232,1,L_SIZE),
				to_sfixed(0.2236,1,L_SIZE),
				to_sfixed(0.2239,1,L_SIZE),
				to_sfixed(0.2243,1,L_SIZE),
				to_sfixed(0.2246,1,L_SIZE),
				to_sfixed(0.2250,1,L_SIZE),
				to_sfixed(0.2253,1,L_SIZE),
				to_sfixed(0.2257,1,L_SIZE),
				to_sfixed(0.2260,1,L_SIZE),
				to_sfixed(0.2264,1,L_SIZE),
				to_sfixed(0.2267,1,L_SIZE),
				to_sfixed(0.2271,1,L_SIZE),
				to_sfixed(0.2274,1,L_SIZE),
				to_sfixed(0.2277,1,L_SIZE),
				to_sfixed(0.2281,1,L_SIZE),
				to_sfixed(0.2284,1,L_SIZE),
				to_sfixed(0.2288,1,L_SIZE),
				to_sfixed(0.2291,1,L_SIZE),
				to_sfixed(0.2295,1,L_SIZE),
				to_sfixed(0.2298,1,L_SIZE),
				to_sfixed(0.2302,1,L_SIZE),
				to_sfixed(0.2305,1,L_SIZE),
				to_sfixed(0.2309,1,L_SIZE),
				to_sfixed(0.2312,1,L_SIZE),
				to_sfixed(0.2316,1,L_SIZE),
				to_sfixed(0.2319,1,L_SIZE),
				to_sfixed(0.2323,1,L_SIZE),
				to_sfixed(0.2326,1,L_SIZE),
				to_sfixed(0.2329,1,L_SIZE),
				to_sfixed(0.2333,1,L_SIZE),
				to_sfixed(0.2336,1,L_SIZE),
				to_sfixed(0.2340,1,L_SIZE),
				to_sfixed(0.2343,1,L_SIZE),
				to_sfixed(0.2347,1,L_SIZE),
				to_sfixed(0.2350,1,L_SIZE),
				to_sfixed(0.2354,1,L_SIZE),
				to_sfixed(0.2357,1,L_SIZE),
				to_sfixed(0.2361,1,L_SIZE),
				to_sfixed(0.2364,1,L_SIZE),
				to_sfixed(0.2368,1,L_SIZE),
				to_sfixed(0.2371,1,L_SIZE),
				to_sfixed(0.2374,1,L_SIZE),
				to_sfixed(0.2378,1,L_SIZE),
				to_sfixed(0.2381,1,L_SIZE),
				to_sfixed(0.2385,1,L_SIZE),
				to_sfixed(0.2388,1,L_SIZE),
				to_sfixed(0.2392,1,L_SIZE),
				to_sfixed(0.2395,1,L_SIZE),
				to_sfixed(0.2399,1,L_SIZE),
				to_sfixed(0.2402,1,L_SIZE),
				to_sfixed(0.2406,1,L_SIZE),
				to_sfixed(0.2409,1,L_SIZE),
				to_sfixed(0.2412,1,L_SIZE),
				to_sfixed(0.2416,1,L_SIZE),
				to_sfixed(0.2419,1,L_SIZE),
				to_sfixed(0.2423,1,L_SIZE),
				to_sfixed(0.2426,1,L_SIZE),
				to_sfixed(0.2430,1,L_SIZE),
				to_sfixed(0.2433,1,L_SIZE),
				to_sfixed(0.2437,1,L_SIZE),
				to_sfixed(0.2440,1,L_SIZE),
				to_sfixed(0.2443,1,L_SIZE),
				to_sfixed(0.2447,1,L_SIZE),
				to_sfixed(0.2450,1,L_SIZE),
				to_sfixed(0.2454,1,L_SIZE),
				to_sfixed(0.2457,1,L_SIZE),
				to_sfixed(0.2461,1,L_SIZE),
				to_sfixed(0.2464,1,L_SIZE),
				to_sfixed(0.2468,1,L_SIZE),
				to_sfixed(0.2471,1,L_SIZE),
				to_sfixed(0.2474,1,L_SIZE),
				to_sfixed(0.2478,1,L_SIZE),
				to_sfixed(0.2481,1,L_SIZE),
				to_sfixed(0.2485,1,L_SIZE),
				to_sfixed(0.2488,1,L_SIZE),
				to_sfixed(0.2492,1,L_SIZE),
				to_sfixed(0.2495,1,L_SIZE),
				to_sfixed(0.2498,1,L_SIZE),
				to_sfixed(0.2502,1,L_SIZE),
				to_sfixed(0.2505,1,L_SIZE),
				to_sfixed(0.2509,1,L_SIZE),
				to_sfixed(0.2512,1,L_SIZE),
				to_sfixed(0.2516,1,L_SIZE),
				to_sfixed(0.2519,1,L_SIZE),
				to_sfixed(0.2522,1,L_SIZE),
				to_sfixed(0.2526,1,L_SIZE),
				to_sfixed(0.2529,1,L_SIZE),
				to_sfixed(0.2533,1,L_SIZE),
				to_sfixed(0.2536,1,L_SIZE),
				to_sfixed(0.2540,1,L_SIZE),
				to_sfixed(0.2543,1,L_SIZE),
				to_sfixed(0.2546,1,L_SIZE),
				to_sfixed(0.2550,1,L_SIZE),
				to_sfixed(0.2553,1,L_SIZE),
				to_sfixed(0.2557,1,L_SIZE),
				to_sfixed(0.2560,1,L_SIZE),
				to_sfixed(0.2564,1,L_SIZE),
				to_sfixed(0.2567,1,L_SIZE),
				to_sfixed(0.2570,1,L_SIZE),
				to_sfixed(0.2574,1,L_SIZE),
				to_sfixed(0.2577,1,L_SIZE),
				to_sfixed(0.2581,1,L_SIZE),
				to_sfixed(0.2584,1,L_SIZE),
				to_sfixed(0.2588,1,L_SIZE),
				to_sfixed(0.2591,1,L_SIZE),
				to_sfixed(0.2594,1,L_SIZE),
				to_sfixed(0.2598,1,L_SIZE),
				to_sfixed(0.2601,1,L_SIZE),
				to_sfixed(0.2605,1,L_SIZE),
				to_sfixed(0.2608,1,L_SIZE),
				to_sfixed(0.2611,1,L_SIZE),
				to_sfixed(0.2615,1,L_SIZE),
				to_sfixed(0.2618,1,L_SIZE),
				to_sfixed(0.2622,1,L_SIZE),
				to_sfixed(0.2625,1,L_SIZE),
				to_sfixed(0.2628,1,L_SIZE),
				to_sfixed(0.2632,1,L_SIZE),
				to_sfixed(0.2635,1,L_SIZE),
				to_sfixed(0.2639,1,L_SIZE),
				to_sfixed(0.2642,1,L_SIZE),
				to_sfixed(0.2646,1,L_SIZE),
				to_sfixed(0.2649,1,L_SIZE),
				to_sfixed(0.2652,1,L_SIZE),
				to_sfixed(0.2656,1,L_SIZE),
				to_sfixed(0.2659,1,L_SIZE),
				to_sfixed(0.2663,1,L_SIZE),
				to_sfixed(0.2666,1,L_SIZE),
				to_sfixed(0.2669,1,L_SIZE),
				to_sfixed(0.2673,1,L_SIZE),
				to_sfixed(0.2676,1,L_SIZE),
				to_sfixed(0.2680,1,L_SIZE),
				to_sfixed(0.2683,1,L_SIZE),
				to_sfixed(0.2686,1,L_SIZE),
				to_sfixed(0.2690,1,L_SIZE),
				to_sfixed(0.2693,1,L_SIZE),
				to_sfixed(0.2697,1,L_SIZE),
				to_sfixed(0.2700,1,L_SIZE),
				to_sfixed(0.2703,1,L_SIZE),
				to_sfixed(0.2707,1,L_SIZE),
				to_sfixed(0.2710,1,L_SIZE),
				to_sfixed(0.2713,1,L_SIZE),
				to_sfixed(0.2717,1,L_SIZE),
				to_sfixed(0.2720,1,L_SIZE),
				to_sfixed(0.2724,1,L_SIZE),
				to_sfixed(0.2727,1,L_SIZE),
				to_sfixed(0.2730,1,L_SIZE),
				to_sfixed(0.2734,1,L_SIZE),
				to_sfixed(0.2737,1,L_SIZE),
				to_sfixed(0.2741,1,L_SIZE),
				to_sfixed(0.2744,1,L_SIZE),
				to_sfixed(0.2747,1,L_SIZE),
				to_sfixed(0.2751,1,L_SIZE),
				to_sfixed(0.2754,1,L_SIZE),
				to_sfixed(0.2758,1,L_SIZE),
				to_sfixed(0.2761,1,L_SIZE),
				to_sfixed(0.2764,1,L_SIZE),
				to_sfixed(0.2768,1,L_SIZE),
				to_sfixed(0.2771,1,L_SIZE),
				to_sfixed(0.2774,1,L_SIZE),
				to_sfixed(0.2778,1,L_SIZE),
				to_sfixed(0.2781,1,L_SIZE),
				to_sfixed(0.2785,1,L_SIZE),
				to_sfixed(0.2788,1,L_SIZE),
				to_sfixed(0.2791,1,L_SIZE),
				to_sfixed(0.2795,1,L_SIZE),
				to_sfixed(0.2798,1,L_SIZE),
				to_sfixed(0.2801,1,L_SIZE),
				to_sfixed(0.2805,1,L_SIZE),
				to_sfixed(0.2808,1,L_SIZE),
				to_sfixed(0.2812,1,L_SIZE),
				to_sfixed(0.2815,1,L_SIZE),
				to_sfixed(0.2818,1,L_SIZE),
				to_sfixed(0.2822,1,L_SIZE),
				to_sfixed(0.2825,1,L_SIZE),
				to_sfixed(0.2828,1,L_SIZE),
				to_sfixed(0.2832,1,L_SIZE),
				to_sfixed(0.2835,1,L_SIZE),
				to_sfixed(0.2839,1,L_SIZE),
				to_sfixed(0.2842,1,L_SIZE),
				to_sfixed(0.2845,1,L_SIZE),
				to_sfixed(0.2849,1,L_SIZE),
				to_sfixed(0.2852,1,L_SIZE),
				to_sfixed(0.2855,1,L_SIZE),
				to_sfixed(0.2859,1,L_SIZE),
				to_sfixed(0.2862,1,L_SIZE),
				to_sfixed(0.2865,1,L_SIZE),
				to_sfixed(0.2869,1,L_SIZE),
				to_sfixed(0.2872,1,L_SIZE),
				to_sfixed(0.2876,1,L_SIZE),
				to_sfixed(0.2879,1,L_SIZE),
				to_sfixed(0.2882,1,L_SIZE),
				to_sfixed(0.2886,1,L_SIZE),
				to_sfixed(0.2889,1,L_SIZE),
				to_sfixed(0.2892,1,L_SIZE),
				to_sfixed(0.2896,1,L_SIZE),
				to_sfixed(0.2899,1,L_SIZE),
				to_sfixed(0.2902,1,L_SIZE),
				to_sfixed(0.2906,1,L_SIZE),
				to_sfixed(0.2909,1,L_SIZE),
				to_sfixed(0.2912,1,L_SIZE),
				to_sfixed(0.2916,1,L_SIZE),
				to_sfixed(0.2919,1,L_SIZE),
				to_sfixed(0.2923,1,L_SIZE),
				to_sfixed(0.2926,1,L_SIZE),
				to_sfixed(0.2929,1,L_SIZE),
				to_sfixed(0.2933,1,L_SIZE),
				to_sfixed(0.2936,1,L_SIZE),
				to_sfixed(0.2939,1,L_SIZE),
				to_sfixed(0.2943,1,L_SIZE),
				to_sfixed(0.2946,1,L_SIZE),
				to_sfixed(0.2949,1,L_SIZE),
				to_sfixed(0.2953,1,L_SIZE),
				to_sfixed(0.2956,1,L_SIZE),
				to_sfixed(0.2959,1,L_SIZE),
				to_sfixed(0.2963,1,L_SIZE),
				to_sfixed(0.2966,1,L_SIZE),
				to_sfixed(0.2969,1,L_SIZE),
				to_sfixed(0.2973,1,L_SIZE),
				to_sfixed(0.2976,1,L_SIZE),
				to_sfixed(0.2979,1,L_SIZE),
				to_sfixed(0.2983,1,L_SIZE),
				to_sfixed(0.2986,1,L_SIZE),
				to_sfixed(0.2989,1,L_SIZE),
				to_sfixed(0.2993,1,L_SIZE),
				to_sfixed(0.2996,1,L_SIZE),
				to_sfixed(0.2999,1,L_SIZE),
				to_sfixed(0.3003,1,L_SIZE),
				to_sfixed(0.3006,1,L_SIZE),
				to_sfixed(0.3009,1,L_SIZE),
				to_sfixed(0.3013,1,L_SIZE),
				to_sfixed(0.3016,1,L_SIZE),
				to_sfixed(0.3019,1,L_SIZE),
				to_sfixed(0.3023,1,L_SIZE),
				to_sfixed(0.3026,1,L_SIZE),
				to_sfixed(0.3029,1,L_SIZE),
				to_sfixed(0.3033,1,L_SIZE),
				to_sfixed(0.3036,1,L_SIZE),
				to_sfixed(0.3039,1,L_SIZE),
				to_sfixed(0.3043,1,L_SIZE),
				to_sfixed(0.3046,1,L_SIZE),
				to_sfixed(0.3049,1,L_SIZE),
				to_sfixed(0.3053,1,L_SIZE),
				to_sfixed(0.3056,1,L_SIZE),
				to_sfixed(0.3059,1,L_SIZE),
				to_sfixed(0.3063,1,L_SIZE),
				to_sfixed(0.3066,1,L_SIZE),
				to_sfixed(0.3069,1,L_SIZE),
				to_sfixed(0.3072,1,L_SIZE),
				to_sfixed(0.3076,1,L_SIZE),
				to_sfixed(0.3079,1,L_SIZE),
				to_sfixed(0.3082,1,L_SIZE),
				to_sfixed(0.3086,1,L_SIZE),
				to_sfixed(0.3089,1,L_SIZE),
				to_sfixed(0.3092,1,L_SIZE),
				to_sfixed(0.3096,1,L_SIZE),
				to_sfixed(0.3099,1,L_SIZE),
				to_sfixed(0.3102,1,L_SIZE),
				to_sfixed(0.3106,1,L_SIZE),
				to_sfixed(0.3109,1,L_SIZE),
				to_sfixed(0.3112,1,L_SIZE),
				to_sfixed(0.3116,1,L_SIZE),
				to_sfixed(0.3119,1,L_SIZE),
				to_sfixed(0.3122,1,L_SIZE),
				to_sfixed(0.3125,1,L_SIZE),
				to_sfixed(0.3129,1,L_SIZE),
				to_sfixed(0.3132,1,L_SIZE),
				to_sfixed(0.3135,1,L_SIZE),
				to_sfixed(0.3139,1,L_SIZE),
				to_sfixed(0.3142,1,L_SIZE),
				to_sfixed(0.3145,1,L_SIZE),
				to_sfixed(0.3149,1,L_SIZE),
				to_sfixed(0.3152,1,L_SIZE),
				to_sfixed(0.3155,1,L_SIZE),
				to_sfixed(0.3158,1,L_SIZE),
				to_sfixed(0.3162,1,L_SIZE),
				to_sfixed(0.3165,1,L_SIZE),
				to_sfixed(0.3168,1,L_SIZE),
				to_sfixed(0.3172,1,L_SIZE),
				to_sfixed(0.3175,1,L_SIZE),
				to_sfixed(0.3178,1,L_SIZE),
				to_sfixed(0.3182,1,L_SIZE),
				to_sfixed(0.3185,1,L_SIZE),
				to_sfixed(0.3188,1,L_SIZE),
				to_sfixed(0.3191,1,L_SIZE),
				to_sfixed(0.3195,1,L_SIZE),
				to_sfixed(0.3198,1,L_SIZE),
				to_sfixed(0.3201,1,L_SIZE),
				to_sfixed(0.3205,1,L_SIZE),
				to_sfixed(0.3208,1,L_SIZE),
				to_sfixed(0.3211,1,L_SIZE),
				to_sfixed(0.3214,1,L_SIZE),
				to_sfixed(0.3218,1,L_SIZE),
				to_sfixed(0.3221,1,L_SIZE),
				to_sfixed(0.3224,1,L_SIZE),
				to_sfixed(0.3228,1,L_SIZE),
				to_sfixed(0.3231,1,L_SIZE),
				to_sfixed(0.3234,1,L_SIZE),
				to_sfixed(0.3237,1,L_SIZE),
				to_sfixed(0.3241,1,L_SIZE),
				to_sfixed(0.3244,1,L_SIZE),
				to_sfixed(0.3247,1,L_SIZE),
				to_sfixed(0.3250,1,L_SIZE),
				to_sfixed(0.3254,1,L_SIZE),
				to_sfixed(0.3257,1,L_SIZE),
				to_sfixed(0.3260,1,L_SIZE),
				to_sfixed(0.3264,1,L_SIZE),
				to_sfixed(0.3267,1,L_SIZE),
				to_sfixed(0.3270,1,L_SIZE),
				to_sfixed(0.3273,1,L_SIZE),
				to_sfixed(0.3277,1,L_SIZE),
				to_sfixed(0.3280,1,L_SIZE),
				to_sfixed(0.3283,1,L_SIZE),
				to_sfixed(0.3286,1,L_SIZE),
				to_sfixed(0.3290,1,L_SIZE),
				to_sfixed(0.3293,1,L_SIZE),
				to_sfixed(0.3296,1,L_SIZE),
				to_sfixed(0.3300,1,L_SIZE),
				to_sfixed(0.3303,1,L_SIZE),
				to_sfixed(0.3306,1,L_SIZE),
				to_sfixed(0.3309,1,L_SIZE),
				to_sfixed(0.3313,1,L_SIZE),
				to_sfixed(0.3316,1,L_SIZE),
				to_sfixed(0.3319,1,L_SIZE),
				to_sfixed(0.3322,1,L_SIZE),
				to_sfixed(0.3326,1,L_SIZE),
				to_sfixed(0.3329,1,L_SIZE),
				to_sfixed(0.3332,1,L_SIZE),
				to_sfixed(0.3335,1,L_SIZE),
				to_sfixed(0.3339,1,L_SIZE),
				to_sfixed(0.3342,1,L_SIZE),
				to_sfixed(0.3345,1,L_SIZE),
				to_sfixed(0.3348,1,L_SIZE),
				to_sfixed(0.3352,1,L_SIZE),
				to_sfixed(0.3355,1,L_SIZE),
				to_sfixed(0.3358,1,L_SIZE),
				to_sfixed(0.3361,1,L_SIZE),
				to_sfixed(0.3365,1,L_SIZE),
				to_sfixed(0.3368,1,L_SIZE),
				to_sfixed(0.3371,1,L_SIZE),
				to_sfixed(0.3374,1,L_SIZE),
				to_sfixed(0.3378,1,L_SIZE),
				to_sfixed(0.3381,1,L_SIZE),
				to_sfixed(0.3384,1,L_SIZE),
				to_sfixed(0.3387,1,L_SIZE),
				to_sfixed(0.3391,1,L_SIZE),
				to_sfixed(0.3394,1,L_SIZE),
				to_sfixed(0.3397,1,L_SIZE),
				to_sfixed(0.3400,1,L_SIZE),
				to_sfixed(0.3404,1,L_SIZE),
				to_sfixed(0.3407,1,L_SIZE),
				to_sfixed(0.3410,1,L_SIZE),
				to_sfixed(0.3413,1,L_SIZE),
				to_sfixed(0.3416,1,L_SIZE),
				to_sfixed(0.3420,1,L_SIZE),
				to_sfixed(0.3423,1,L_SIZE),
				to_sfixed(0.3426,1,L_SIZE),
				to_sfixed(0.3429,1,L_SIZE),
				to_sfixed(0.3433,1,L_SIZE),
				to_sfixed(0.3436,1,L_SIZE),
				to_sfixed(0.3439,1,L_SIZE),
				to_sfixed(0.3442,1,L_SIZE),
				to_sfixed(0.3446,1,L_SIZE),
				to_sfixed(0.3449,1,L_SIZE),
				to_sfixed(0.3452,1,L_SIZE),
				to_sfixed(0.3455,1,L_SIZE),
				to_sfixed(0.3458,1,L_SIZE),
				to_sfixed(0.3462,1,L_SIZE),
				to_sfixed(0.3465,1,L_SIZE),
				to_sfixed(0.3468,1,L_SIZE),
				to_sfixed(0.3471,1,L_SIZE),
				to_sfixed(0.3475,1,L_SIZE),
				to_sfixed(0.3478,1,L_SIZE),
				to_sfixed(0.3481,1,L_SIZE),
				to_sfixed(0.3484,1,L_SIZE),
				to_sfixed(0.3487,1,L_SIZE),
				to_sfixed(0.3491,1,L_SIZE),
				to_sfixed(0.3494,1,L_SIZE),
				to_sfixed(0.3497,1,L_SIZE),
				to_sfixed(0.3500,1,L_SIZE),
				to_sfixed(0.3504,1,L_SIZE),
				to_sfixed(0.3507,1,L_SIZE),
				to_sfixed(0.3510,1,L_SIZE),
				to_sfixed(0.3513,1,L_SIZE),
				to_sfixed(0.3516,1,L_SIZE),
				to_sfixed(0.3520,1,L_SIZE),
				to_sfixed(0.3523,1,L_SIZE),
				to_sfixed(0.3526,1,L_SIZE),
				to_sfixed(0.3529,1,L_SIZE),
				to_sfixed(0.3532,1,L_SIZE),
				to_sfixed(0.3536,1,L_SIZE),
				to_sfixed(0.3539,1,L_SIZE),
				to_sfixed(0.3542,1,L_SIZE),
				to_sfixed(0.3545,1,L_SIZE),
				to_sfixed(0.3548,1,L_SIZE),
				to_sfixed(0.3552,1,L_SIZE),
				to_sfixed(0.3555,1,L_SIZE),
				to_sfixed(0.3558,1,L_SIZE),
				to_sfixed(0.3561,1,L_SIZE),
				to_sfixed(0.3564,1,L_SIZE),
				to_sfixed(0.3568,1,L_SIZE),
				to_sfixed(0.3571,1,L_SIZE),
				to_sfixed(0.3574,1,L_SIZE),
				to_sfixed(0.3577,1,L_SIZE),
				to_sfixed(0.3580,1,L_SIZE),
				to_sfixed(0.3584,1,L_SIZE),
				to_sfixed(0.3587,1,L_SIZE),
				to_sfixed(0.3590,1,L_SIZE),
				to_sfixed(0.3593,1,L_SIZE),
				to_sfixed(0.3596,1,L_SIZE),
				to_sfixed(0.3600,1,L_SIZE),
				to_sfixed(0.3603,1,L_SIZE),
				to_sfixed(0.3606,1,L_SIZE),
				to_sfixed(0.3609,1,L_SIZE),
				to_sfixed(0.3612,1,L_SIZE),
				to_sfixed(0.3615,1,L_SIZE),
				to_sfixed(0.3619,1,L_SIZE),
				to_sfixed(0.3622,1,L_SIZE),
				to_sfixed(0.3625,1,L_SIZE),
				to_sfixed(0.3628,1,L_SIZE),
				to_sfixed(0.3631,1,L_SIZE),
				to_sfixed(0.3635,1,L_SIZE),
				to_sfixed(0.3638,1,L_SIZE),
				to_sfixed(0.3641,1,L_SIZE),
				to_sfixed(0.3644,1,L_SIZE),
				to_sfixed(0.3647,1,L_SIZE),
				to_sfixed(0.3650,1,L_SIZE),
				to_sfixed(0.3654,1,L_SIZE),
				to_sfixed(0.3657,1,L_SIZE),
				to_sfixed(0.3660,1,L_SIZE),
				to_sfixed(0.3663,1,L_SIZE),
				to_sfixed(0.3666,1,L_SIZE),
				to_sfixed(0.3669,1,L_SIZE),
				to_sfixed(0.3673,1,L_SIZE),
				to_sfixed(0.3676,1,L_SIZE),
				to_sfixed(0.3679,1,L_SIZE),
				to_sfixed(0.3682,1,L_SIZE),
				to_sfixed(0.3685,1,L_SIZE),
				to_sfixed(0.3688,1,L_SIZE),
				to_sfixed(0.3692,1,L_SIZE),
				to_sfixed(0.3695,1,L_SIZE),
				to_sfixed(0.3698,1,L_SIZE),
				to_sfixed(0.3701,1,L_SIZE),
				to_sfixed(0.3704,1,L_SIZE),
				to_sfixed(0.3707,1,L_SIZE),
				to_sfixed(0.3711,1,L_SIZE),
				to_sfixed(0.3714,1,L_SIZE),
				to_sfixed(0.3717,1,L_SIZE),
				to_sfixed(0.3720,1,L_SIZE),
				to_sfixed(0.3723,1,L_SIZE),
				to_sfixed(0.3726,1,L_SIZE),
				to_sfixed(0.3730,1,L_SIZE),
				to_sfixed(0.3733,1,L_SIZE),
				to_sfixed(0.3736,1,L_SIZE),
				to_sfixed(0.3739,1,L_SIZE),
				to_sfixed(0.3742,1,L_SIZE),
				to_sfixed(0.3745,1,L_SIZE),
				to_sfixed(0.3748,1,L_SIZE),
				to_sfixed(0.3752,1,L_SIZE),
				to_sfixed(0.3755,1,L_SIZE),
				to_sfixed(0.3758,1,L_SIZE),
				to_sfixed(0.3761,1,L_SIZE),
				to_sfixed(0.3764,1,L_SIZE),
				to_sfixed(0.3767,1,L_SIZE),
				to_sfixed(0.3770,1,L_SIZE),
				to_sfixed(0.3774,1,L_SIZE),
				to_sfixed(0.3777,1,L_SIZE),
				to_sfixed(0.3780,1,L_SIZE),
				to_sfixed(0.3783,1,L_SIZE),
				to_sfixed(0.3786,1,L_SIZE),
				to_sfixed(0.3789,1,L_SIZE),
				to_sfixed(0.3792,1,L_SIZE),
				to_sfixed(0.3796,1,L_SIZE),
				to_sfixed(0.3799,1,L_SIZE),
				to_sfixed(0.3802,1,L_SIZE),
				to_sfixed(0.3805,1,L_SIZE),
				to_sfixed(0.3808,1,L_SIZE),
				to_sfixed(0.3811,1,L_SIZE),
				to_sfixed(0.3814,1,L_SIZE),
				to_sfixed(0.3817,1,L_SIZE),
				to_sfixed(0.3821,1,L_SIZE),
				to_sfixed(0.3824,1,L_SIZE),
				to_sfixed(0.3827,1,L_SIZE),
				to_sfixed(0.3830,1,L_SIZE),
				to_sfixed(0.3833,1,L_SIZE),
				to_sfixed(0.3836,1,L_SIZE),
				to_sfixed(0.3839,1,L_SIZE),
				to_sfixed(0.3842,1,L_SIZE),
				to_sfixed(0.3846,1,L_SIZE),
				to_sfixed(0.3849,1,L_SIZE),
				to_sfixed(0.3852,1,L_SIZE),
				to_sfixed(0.3855,1,L_SIZE),
				to_sfixed(0.3858,1,L_SIZE),
				to_sfixed(0.3861,1,L_SIZE),
				to_sfixed(0.3864,1,L_SIZE),
				to_sfixed(0.3867,1,L_SIZE),
				to_sfixed(0.3870,1,L_SIZE),
				to_sfixed(0.3874,1,L_SIZE),
				to_sfixed(0.3877,1,L_SIZE),
				to_sfixed(0.3880,1,L_SIZE),
				to_sfixed(0.3883,1,L_SIZE),
				to_sfixed(0.3886,1,L_SIZE),
				to_sfixed(0.3889,1,L_SIZE),
				to_sfixed(0.3892,1,L_SIZE),
				to_sfixed(0.3895,1,L_SIZE),
				to_sfixed(0.3898,1,L_SIZE),
				to_sfixed(0.3902,1,L_SIZE),
				to_sfixed(0.3905,1,L_SIZE),
				to_sfixed(0.3908,1,L_SIZE),
				to_sfixed(0.3911,1,L_SIZE),
				to_sfixed(0.3914,1,L_SIZE),
				to_sfixed(0.3917,1,L_SIZE),
				to_sfixed(0.3920,1,L_SIZE),
				to_sfixed(0.3923,1,L_SIZE),
				to_sfixed(0.3926,1,L_SIZE),
				to_sfixed(0.3929,1,L_SIZE),
				to_sfixed(0.3933,1,L_SIZE),
				to_sfixed(0.3936,1,L_SIZE),
				to_sfixed(0.3939,1,L_SIZE),
				to_sfixed(0.3942,1,L_SIZE),
				to_sfixed(0.3945,1,L_SIZE),
				to_sfixed(0.3948,1,L_SIZE),
				to_sfixed(0.3951,1,L_SIZE),
				to_sfixed(0.3954,1,L_SIZE),
				to_sfixed(0.3957,1,L_SIZE),
				to_sfixed(0.3960,1,L_SIZE),
				to_sfixed(0.3964,1,L_SIZE),
				to_sfixed(0.3967,1,L_SIZE),
				to_sfixed(0.3970,1,L_SIZE),
				to_sfixed(0.3973,1,L_SIZE),
				to_sfixed(0.3976,1,L_SIZE),
				to_sfixed(0.3979,1,L_SIZE),
				to_sfixed(0.3982,1,L_SIZE),
				to_sfixed(0.3985,1,L_SIZE),
				to_sfixed(0.3988,1,L_SIZE),
				to_sfixed(0.3991,1,L_SIZE),
				to_sfixed(0.3994,1,L_SIZE),
				to_sfixed(0.3997,1,L_SIZE),
				to_sfixed(0.4000,1,L_SIZE),
				to_sfixed(0.4004,1,L_SIZE),
				to_sfixed(0.4007,1,L_SIZE),
				to_sfixed(0.4010,1,L_SIZE),
				to_sfixed(0.4013,1,L_SIZE),
				to_sfixed(0.4016,1,L_SIZE),
				to_sfixed(0.4019,1,L_SIZE),
				to_sfixed(0.4022,1,L_SIZE),
				to_sfixed(0.4025,1,L_SIZE),
				to_sfixed(0.4028,1,L_SIZE),
				to_sfixed(0.4031,1,L_SIZE),
				to_sfixed(0.4034,1,L_SIZE),
				to_sfixed(0.4037,1,L_SIZE),
				to_sfixed(0.4040,1,L_SIZE),
				to_sfixed(0.4043,1,L_SIZE),
				to_sfixed(0.4047,1,L_SIZE),
				to_sfixed(0.4050,1,L_SIZE),
				to_sfixed(0.4053,1,L_SIZE),
				to_sfixed(0.4056,1,L_SIZE),
				to_sfixed(0.4059,1,L_SIZE),
				to_sfixed(0.4062,1,L_SIZE),
				to_sfixed(0.4065,1,L_SIZE),
				to_sfixed(0.4068,1,L_SIZE),
				to_sfixed(0.4071,1,L_SIZE),
				to_sfixed(0.4074,1,L_SIZE),
				to_sfixed(0.4077,1,L_SIZE),
				to_sfixed(0.4080,1,L_SIZE),
				to_sfixed(0.4083,1,L_SIZE),
				to_sfixed(0.4086,1,L_SIZE),
				to_sfixed(0.4089,1,L_SIZE),
				to_sfixed(0.4092,1,L_SIZE),
				to_sfixed(0.4095,1,L_SIZE),
				to_sfixed(0.4098,1,L_SIZE),
				to_sfixed(0.4101,1,L_SIZE),
				to_sfixed(0.4105,1,L_SIZE),
				to_sfixed(0.4108,1,L_SIZE),
				to_sfixed(0.4111,1,L_SIZE),
				to_sfixed(0.4114,1,L_SIZE),
				to_sfixed(0.4117,1,L_SIZE),
				to_sfixed(0.4120,1,L_SIZE),
				to_sfixed(0.4123,1,L_SIZE),
				to_sfixed(0.4126,1,L_SIZE),
				to_sfixed(0.4129,1,L_SIZE),
				to_sfixed(0.4132,1,L_SIZE),
				to_sfixed(0.4135,1,L_SIZE),
				to_sfixed(0.4138,1,L_SIZE),
				to_sfixed(0.4141,1,L_SIZE),
				to_sfixed(0.4144,1,L_SIZE),
				to_sfixed(0.4147,1,L_SIZE),
				to_sfixed(0.4150,1,L_SIZE),
				to_sfixed(0.4153,1,L_SIZE),
				to_sfixed(0.4156,1,L_SIZE),
				to_sfixed(0.4159,1,L_SIZE),
				to_sfixed(0.4162,1,L_SIZE),
				to_sfixed(0.4165,1,L_SIZE),
				to_sfixed(0.4168,1,L_SIZE),
				to_sfixed(0.4171,1,L_SIZE),
				to_sfixed(0.4174,1,L_SIZE),
				to_sfixed(0.4177,1,L_SIZE),
				to_sfixed(0.4180,1,L_SIZE),
				to_sfixed(0.4183,1,L_SIZE),
				to_sfixed(0.4186,1,L_SIZE),
				to_sfixed(0.4189,1,L_SIZE),
				to_sfixed(0.4192,1,L_SIZE),
				to_sfixed(0.4195,1,L_SIZE),
				to_sfixed(0.4198,1,L_SIZE),
				to_sfixed(0.4202,1,L_SIZE),
				to_sfixed(0.4205,1,L_SIZE),
				to_sfixed(0.4208,1,L_SIZE),
				to_sfixed(0.4211,1,L_SIZE),
				to_sfixed(0.4214,1,L_SIZE),
				to_sfixed(0.4217,1,L_SIZE),
				to_sfixed(0.4220,1,L_SIZE),
				to_sfixed(0.4223,1,L_SIZE),
				to_sfixed(0.4226,1,L_SIZE),
				to_sfixed(0.4229,1,L_SIZE),
				to_sfixed(0.4232,1,L_SIZE),
				to_sfixed(0.4235,1,L_SIZE),
				to_sfixed(0.4238,1,L_SIZE),
				to_sfixed(0.4241,1,L_SIZE),
				to_sfixed(0.4244,1,L_SIZE),
				to_sfixed(0.4247,1,L_SIZE),
				to_sfixed(0.4250,1,L_SIZE),
				to_sfixed(0.4253,1,L_SIZE),
				to_sfixed(0.4256,1,L_SIZE),
				to_sfixed(0.4259,1,L_SIZE),
				to_sfixed(0.4262,1,L_SIZE),
				to_sfixed(0.4265,1,L_SIZE),
				to_sfixed(0.4268,1,L_SIZE),
				to_sfixed(0.4271,1,L_SIZE),
				to_sfixed(0.4274,1,L_SIZE),
				to_sfixed(0.4277,1,L_SIZE),
				to_sfixed(0.4280,1,L_SIZE),
				to_sfixed(0.4283,1,L_SIZE),
				to_sfixed(0.4286,1,L_SIZE),
				to_sfixed(0.4289,1,L_SIZE),
				to_sfixed(0.4292,1,L_SIZE),
				to_sfixed(0.4295,1,L_SIZE),
				to_sfixed(0.4298,1,L_SIZE),
				to_sfixed(0.4301,1,L_SIZE),
				to_sfixed(0.4304,1,L_SIZE),
				to_sfixed(0.4306,1,L_SIZE),
				to_sfixed(0.4309,1,L_SIZE),
				to_sfixed(0.4312,1,L_SIZE),
				to_sfixed(0.4315,1,L_SIZE),
				to_sfixed(0.4318,1,L_SIZE),
				to_sfixed(0.4321,1,L_SIZE),
				to_sfixed(0.4324,1,L_SIZE),
				to_sfixed(0.4327,1,L_SIZE),
				to_sfixed(0.4330,1,L_SIZE),
				to_sfixed(0.4333,1,L_SIZE),
				to_sfixed(0.4336,1,L_SIZE),
				to_sfixed(0.4339,1,L_SIZE),
				to_sfixed(0.4342,1,L_SIZE),
				to_sfixed(0.4345,1,L_SIZE),
				to_sfixed(0.4348,1,L_SIZE),
				to_sfixed(0.4351,1,L_SIZE),
				to_sfixed(0.4354,1,L_SIZE),
				to_sfixed(0.4357,1,L_SIZE),
				to_sfixed(0.4360,1,L_SIZE),
				to_sfixed(0.4363,1,L_SIZE),
				to_sfixed(0.4366,1,L_SIZE),
				to_sfixed(0.4369,1,L_SIZE),
				to_sfixed(0.4372,1,L_SIZE),
				to_sfixed(0.4375,1,L_SIZE),
				to_sfixed(0.4378,1,L_SIZE),
				to_sfixed(0.4381,1,L_SIZE),
				to_sfixed(0.4384,1,L_SIZE),
				to_sfixed(0.4387,1,L_SIZE),
				to_sfixed(0.4390,1,L_SIZE),
				to_sfixed(0.4393,1,L_SIZE),
				to_sfixed(0.4396,1,L_SIZE),
				to_sfixed(0.4399,1,L_SIZE),
				to_sfixed(0.4401,1,L_SIZE),
				to_sfixed(0.4404,1,L_SIZE),
				to_sfixed(0.4407,1,L_SIZE),
				to_sfixed(0.4410,1,L_SIZE),
				to_sfixed(0.4413,1,L_SIZE),
				to_sfixed(0.4416,1,L_SIZE),
				to_sfixed(0.4419,1,L_SIZE),
				to_sfixed(0.4422,1,L_SIZE),
				to_sfixed(0.4425,1,L_SIZE),
				to_sfixed(0.4428,1,L_SIZE),
				to_sfixed(0.4431,1,L_SIZE),
				to_sfixed(0.4434,1,L_SIZE),
				to_sfixed(0.4437,1,L_SIZE),
				to_sfixed(0.4440,1,L_SIZE),
				to_sfixed(0.4443,1,L_SIZE),
				to_sfixed(0.4446,1,L_SIZE),
				to_sfixed(0.4449,1,L_SIZE),
				to_sfixed(0.4452,1,L_SIZE),
				to_sfixed(0.4454,1,L_SIZE),
				to_sfixed(0.4457,1,L_SIZE),
				to_sfixed(0.4460,1,L_SIZE),
				to_sfixed(0.4463,1,L_SIZE),
				to_sfixed(0.4466,1,L_SIZE),
				to_sfixed(0.4469,1,L_SIZE),
				to_sfixed(0.4472,1,L_SIZE),
				to_sfixed(0.4475,1,L_SIZE),
				to_sfixed(0.4478,1,L_SIZE),
				to_sfixed(0.4481,1,L_SIZE),
				to_sfixed(0.4484,1,L_SIZE),
				to_sfixed(0.4487,1,L_SIZE),
				to_sfixed(0.4490,1,L_SIZE),
				to_sfixed(0.4493,1,L_SIZE),
				to_sfixed(0.4495,1,L_SIZE),
				to_sfixed(0.4498,1,L_SIZE),
				to_sfixed(0.4501,1,L_SIZE),
				to_sfixed(0.4504,1,L_SIZE),
				to_sfixed(0.4507,1,L_SIZE),
				to_sfixed(0.4510,1,L_SIZE),
				to_sfixed(0.4513,1,L_SIZE),
				to_sfixed(0.4516,1,L_SIZE),
				to_sfixed(0.4519,1,L_SIZE),
				to_sfixed(0.4522,1,L_SIZE),
				to_sfixed(0.4525,1,L_SIZE),
				to_sfixed(0.4528,1,L_SIZE),
				to_sfixed(0.4530,1,L_SIZE),
				to_sfixed(0.4533,1,L_SIZE),
				to_sfixed(0.4536,1,L_SIZE),
				to_sfixed(0.4539,1,L_SIZE),
				to_sfixed(0.4542,1,L_SIZE),
				to_sfixed(0.4545,1,L_SIZE),
				to_sfixed(0.4548,1,L_SIZE),
				to_sfixed(0.4551,1,L_SIZE),
				to_sfixed(0.4554,1,L_SIZE),
				to_sfixed(0.4557,1,L_SIZE),
				to_sfixed(0.4560,1,L_SIZE),
				to_sfixed(0.4562,1,L_SIZE),
				to_sfixed(0.4565,1,L_SIZE),
				to_sfixed(0.4568,1,L_SIZE),
				to_sfixed(0.4571,1,L_SIZE),
				to_sfixed(0.4574,1,L_SIZE),
				to_sfixed(0.4577,1,L_SIZE),
				to_sfixed(0.4580,1,L_SIZE),
				to_sfixed(0.4583,1,L_SIZE),
				to_sfixed(0.4586,1,L_SIZE),
				to_sfixed(0.4588,1,L_SIZE),
				to_sfixed(0.4591,1,L_SIZE),
				to_sfixed(0.4594,1,L_SIZE),
				to_sfixed(0.4597,1,L_SIZE),
				to_sfixed(0.4600,1,L_SIZE),
				to_sfixed(0.4603,1,L_SIZE),
				to_sfixed(0.4606,1,L_SIZE),
				to_sfixed(0.4609,1,L_SIZE),
				to_sfixed(0.4612,1,L_SIZE),
				to_sfixed(0.4614,1,L_SIZE),
				to_sfixed(0.4617,1,L_SIZE),
				to_sfixed(0.4620,1,L_SIZE),
				to_sfixed(0.4623,1,L_SIZE),
				to_sfixed(0.4626,1,L_SIZE),
				to_sfixed(0.4629,1,L_SIZE),
				to_sfixed(0.4632,1,L_SIZE),
				to_sfixed(0.4635,1,L_SIZE),
				to_sfixed(0.4637,1,L_SIZE),
				to_sfixed(0.4640,1,L_SIZE),
				to_sfixed(0.4643,1,L_SIZE),
				to_sfixed(0.4646,1,L_SIZE),
				to_sfixed(0.4649,1,L_SIZE),
				to_sfixed(0.4652,1,L_SIZE),
				to_sfixed(0.4655,1,L_SIZE),
				to_sfixed(0.4658,1,L_SIZE),
				to_sfixed(0.4660,1,L_SIZE),
				to_sfixed(0.4663,1,L_SIZE),
				to_sfixed(0.4666,1,L_SIZE),
				to_sfixed(0.4669,1,L_SIZE),
				to_sfixed(0.4672,1,L_SIZE),
				to_sfixed(0.4675,1,L_SIZE),
				to_sfixed(0.4678,1,L_SIZE),
				to_sfixed(0.4680,1,L_SIZE),
				to_sfixed(0.4683,1,L_SIZE),
				to_sfixed(0.4686,1,L_SIZE),
				to_sfixed(0.4689,1,L_SIZE),
				to_sfixed(0.4692,1,L_SIZE),
				to_sfixed(0.4695,1,L_SIZE),
				to_sfixed(0.4698,1,L_SIZE),
				to_sfixed(0.4700,1,L_SIZE),
				to_sfixed(0.4703,1,L_SIZE),
				to_sfixed(0.4706,1,L_SIZE),
				to_sfixed(0.4709,1,L_SIZE),
				to_sfixed(0.4712,1,L_SIZE),
				to_sfixed(0.4715,1,L_SIZE),
				to_sfixed(0.4718,1,L_SIZE),
				to_sfixed(0.4720,1,L_SIZE),
				to_sfixed(0.4723,1,L_SIZE),
				to_sfixed(0.4726,1,L_SIZE),
				to_sfixed(0.4729,1,L_SIZE),
				to_sfixed(0.4732,1,L_SIZE),
				to_sfixed(0.4735,1,L_SIZE),
				to_sfixed(0.4737,1,L_SIZE),
				to_sfixed(0.4740,1,L_SIZE),
				to_sfixed(0.4743,1,L_SIZE),
				to_sfixed(0.4746,1,L_SIZE),
				to_sfixed(0.4749,1,L_SIZE),
				to_sfixed(0.4752,1,L_SIZE),
				to_sfixed(0.4755,1,L_SIZE),
				to_sfixed(0.4757,1,L_SIZE),
				to_sfixed(0.4760,1,L_SIZE),
				to_sfixed(0.4763,1,L_SIZE),
				to_sfixed(0.4766,1,L_SIZE),
				to_sfixed(0.4769,1,L_SIZE),
				to_sfixed(0.4771,1,L_SIZE),
				to_sfixed(0.4774,1,L_SIZE),
				to_sfixed(0.4777,1,L_SIZE),
				to_sfixed(0.4780,1,L_SIZE),
				to_sfixed(0.4783,1,L_SIZE),
				to_sfixed(0.4786,1,L_SIZE),
				to_sfixed(0.4788,1,L_SIZE),
				to_sfixed(0.4791,1,L_SIZE),
				to_sfixed(0.4794,1,L_SIZE),
				to_sfixed(0.4797,1,L_SIZE),
				to_sfixed(0.4800,1,L_SIZE),
				to_sfixed(0.4803,1,L_SIZE),
				to_sfixed(0.4805,1,L_SIZE),
				to_sfixed(0.4808,1,L_SIZE),
				to_sfixed(0.4811,1,L_SIZE),
				to_sfixed(0.4814,1,L_SIZE),
				to_sfixed(0.4817,1,L_SIZE),
				to_sfixed(0.4819,1,L_SIZE),
				to_sfixed(0.4822,1,L_SIZE),
				to_sfixed(0.4825,1,L_SIZE),
				to_sfixed(0.4828,1,L_SIZE),
				to_sfixed(0.4831,1,L_SIZE),
				to_sfixed(0.4833,1,L_SIZE),
				to_sfixed(0.4836,1,L_SIZE),
				to_sfixed(0.4839,1,L_SIZE),
				to_sfixed(0.4842,1,L_SIZE),
				to_sfixed(0.4845,1,L_SIZE),
				to_sfixed(0.4848,1,L_SIZE),
				to_sfixed(0.4850,1,L_SIZE),
				to_sfixed(0.4853,1,L_SIZE),
				to_sfixed(0.4856,1,L_SIZE),
				to_sfixed(0.4859,1,L_SIZE),
				to_sfixed(0.4861,1,L_SIZE),
				to_sfixed(0.4864,1,L_SIZE),
				to_sfixed(0.4867,1,L_SIZE),
				to_sfixed(0.4870,1,L_SIZE),
				to_sfixed(0.4873,1,L_SIZE),
				to_sfixed(0.4875,1,L_SIZE),
				to_sfixed(0.4878,1,L_SIZE),
				to_sfixed(0.4881,1,L_SIZE),
				to_sfixed(0.4884,1,L_SIZE),
				to_sfixed(0.4887,1,L_SIZE),
				to_sfixed(0.4889,1,L_SIZE),
				to_sfixed(0.4892,1,L_SIZE),
				to_sfixed(0.4895,1,L_SIZE),
				to_sfixed(0.4898,1,L_SIZE),
				to_sfixed(0.4901,1,L_SIZE),
				to_sfixed(0.4903,1,L_SIZE),
				to_sfixed(0.4906,1,L_SIZE),
				to_sfixed(0.4909,1,L_SIZE),
				to_sfixed(0.4912,1,L_SIZE),
				to_sfixed(0.4914,1,L_SIZE),
				to_sfixed(0.4917,1,L_SIZE),
				to_sfixed(0.4920,1,L_SIZE),
				to_sfixed(0.4923,1,L_SIZE),
				to_sfixed(0.4926,1,L_SIZE),
				to_sfixed(0.4928,1,L_SIZE),
				to_sfixed(0.4931,1,L_SIZE),
				to_sfixed(0.4934,1,L_SIZE),
				to_sfixed(0.4937,1,L_SIZE),
				to_sfixed(0.4939,1,L_SIZE),
				to_sfixed(0.4942,1,L_SIZE),
				to_sfixed(0.4945,1,L_SIZE),
				to_sfixed(0.4948,1,L_SIZE),
				to_sfixed(0.4950,1,L_SIZE),
				to_sfixed(0.4953,1,L_SIZE),
				to_sfixed(0.4956,1,L_SIZE),
				to_sfixed(0.4959,1,L_SIZE),
				to_sfixed(0.4962,1,L_SIZE),
				to_sfixed(0.4964,1,L_SIZE),
				to_sfixed(0.4967,1,L_SIZE),
				to_sfixed(0.4970,1,L_SIZE),
				to_sfixed(0.4973,1,L_SIZE),
				to_sfixed(0.4975,1,L_SIZE),
				to_sfixed(0.4978,1,L_SIZE),
				to_sfixed(0.4981,1,L_SIZE),
				to_sfixed(0.4984,1,L_SIZE),
				to_sfixed(0.4986,1,L_SIZE),
				to_sfixed(0.4989,1,L_SIZE),
				to_sfixed(0.4992,1,L_SIZE),
				to_sfixed(0.4995,1,L_SIZE),
				to_sfixed(0.4997,1,L_SIZE),
				to_sfixed(0.5000,1,L_SIZE),
				to_sfixed(0.5003,1,L_SIZE),
				to_sfixed(0.5006,1,L_SIZE),
				to_sfixed(0.5008,1,L_SIZE),
				to_sfixed(0.5011,1,L_SIZE),
				to_sfixed(0.5014,1,L_SIZE),
				to_sfixed(0.5017,1,L_SIZE),
				to_sfixed(0.5019,1,L_SIZE),
				to_sfixed(0.5022,1,L_SIZE),
				to_sfixed(0.5025,1,L_SIZE),
				to_sfixed(0.5027,1,L_SIZE),
				to_sfixed(0.5030,1,L_SIZE),
				to_sfixed(0.5033,1,L_SIZE),
				to_sfixed(0.5036,1,L_SIZE),
				to_sfixed(0.5038,1,L_SIZE),
				to_sfixed(0.5041,1,L_SIZE),
				to_sfixed(0.5044,1,L_SIZE),
				to_sfixed(0.5047,1,L_SIZE),
				to_sfixed(0.5049,1,L_SIZE),
				to_sfixed(0.5052,1,L_SIZE),
				to_sfixed(0.5055,1,L_SIZE),
				to_sfixed(0.5058,1,L_SIZE),
				to_sfixed(0.5060,1,L_SIZE),
				to_sfixed(0.5063,1,L_SIZE),
				to_sfixed(0.5066,1,L_SIZE),
				to_sfixed(0.5068,1,L_SIZE),
				to_sfixed(0.5071,1,L_SIZE),
				to_sfixed(0.5074,1,L_SIZE),
				to_sfixed(0.5077,1,L_SIZE),
				to_sfixed(0.5079,1,L_SIZE),
				to_sfixed(0.5082,1,L_SIZE),
				to_sfixed(0.5085,1,L_SIZE),
				to_sfixed(0.5087,1,L_SIZE),
				to_sfixed(0.5090,1,L_SIZE),
				to_sfixed(0.5093,1,L_SIZE),
				to_sfixed(0.5096,1,L_SIZE),
				to_sfixed(0.5098,1,L_SIZE),
				to_sfixed(0.5101,1,L_SIZE),
				to_sfixed(0.5104,1,L_SIZE),
				to_sfixed(0.5106,1,L_SIZE),
				to_sfixed(0.5109,1,L_SIZE),
				to_sfixed(0.5112,1,L_SIZE),
				to_sfixed(0.5115,1,L_SIZE),
				to_sfixed(0.5117,1,L_SIZE),
				to_sfixed(0.5120,1,L_SIZE),
				to_sfixed(0.5123,1,L_SIZE),
				to_sfixed(0.5125,1,L_SIZE),
				to_sfixed(0.5128,1,L_SIZE),
				to_sfixed(0.5131,1,L_SIZE),
				to_sfixed(0.5133,1,L_SIZE),
				to_sfixed(0.5136,1,L_SIZE),
				to_sfixed(0.5139,1,L_SIZE),
				to_sfixed(0.5142,1,L_SIZE),
				to_sfixed(0.5144,1,L_SIZE),
				to_sfixed(0.5147,1,L_SIZE),
				to_sfixed(0.5150,1,L_SIZE),
				to_sfixed(0.5152,1,L_SIZE),
				to_sfixed(0.5155,1,L_SIZE),
				to_sfixed(0.5158,1,L_SIZE),
				to_sfixed(0.5160,1,L_SIZE),
				to_sfixed(0.5163,1,L_SIZE),
				to_sfixed(0.5166,1,L_SIZE),
				to_sfixed(0.5168,1,L_SIZE),
				to_sfixed(0.5171,1,L_SIZE),
				to_sfixed(0.5174,1,L_SIZE),
				to_sfixed(0.5176,1,L_SIZE),
				to_sfixed(0.5179,1,L_SIZE),
				to_sfixed(0.5182,1,L_SIZE),
				to_sfixed(0.5185,1,L_SIZE),
				to_sfixed(0.5187,1,L_SIZE),
				to_sfixed(0.5190,1,L_SIZE),
				to_sfixed(0.5193,1,L_SIZE),
				to_sfixed(0.5195,1,L_SIZE),
				to_sfixed(0.5198,1,L_SIZE),
				to_sfixed(0.5201,1,L_SIZE),
				to_sfixed(0.5203,1,L_SIZE),
				to_sfixed(0.5206,1,L_SIZE),
				to_sfixed(0.5209,1,L_SIZE),
				to_sfixed(0.5211,1,L_SIZE),
				to_sfixed(0.5214,1,L_SIZE),
				to_sfixed(0.5217,1,L_SIZE),
				to_sfixed(0.5219,1,L_SIZE),
				to_sfixed(0.5222,1,L_SIZE),
				to_sfixed(0.5225,1,L_SIZE),
				to_sfixed(0.5227,1,L_SIZE),
				to_sfixed(0.5230,1,L_SIZE),
				to_sfixed(0.5233,1,L_SIZE),
				to_sfixed(0.5235,1,L_SIZE),
				to_sfixed(0.5238,1,L_SIZE),
				to_sfixed(0.5241,1,L_SIZE),
				to_sfixed(0.5243,1,L_SIZE),
				to_sfixed(0.5246,1,L_SIZE),
				to_sfixed(0.5248,1,L_SIZE),
				to_sfixed(0.5251,1,L_SIZE),
				to_sfixed(0.5254,1,L_SIZE),
				to_sfixed(0.5256,1,L_SIZE),
				to_sfixed(0.5259,1,L_SIZE),
				to_sfixed(0.5262,1,L_SIZE),
				to_sfixed(0.5264,1,L_SIZE),
				to_sfixed(0.5267,1,L_SIZE),
				to_sfixed(0.5270,1,L_SIZE),
				to_sfixed(0.5272,1,L_SIZE),
				to_sfixed(0.5275,1,L_SIZE),
				to_sfixed(0.5278,1,L_SIZE),
				to_sfixed(0.5280,1,L_SIZE),
				to_sfixed(0.5283,1,L_SIZE),
				to_sfixed(0.5286,1,L_SIZE),
				to_sfixed(0.5288,1,L_SIZE),
				to_sfixed(0.5291,1,L_SIZE),
				to_sfixed(0.5293,1,L_SIZE),
				to_sfixed(0.5296,1,L_SIZE),
				to_sfixed(0.5299,1,L_SIZE),
				to_sfixed(0.5301,1,L_SIZE),
				to_sfixed(0.5304,1,L_SIZE),
				to_sfixed(0.5307,1,L_SIZE),
				to_sfixed(0.5309,1,L_SIZE),
				to_sfixed(0.5312,1,L_SIZE),
				to_sfixed(0.5314,1,L_SIZE),
				to_sfixed(0.5317,1,L_SIZE),
				to_sfixed(0.5320,1,L_SIZE),
				to_sfixed(0.5322,1,L_SIZE),
				to_sfixed(0.5325,1,L_SIZE),
				to_sfixed(0.5328,1,L_SIZE),
				to_sfixed(0.5330,1,L_SIZE),
				to_sfixed(0.5333,1,L_SIZE),
				to_sfixed(0.5335,1,L_SIZE),
				to_sfixed(0.5338,1,L_SIZE),
				to_sfixed(0.5341,1,L_SIZE),
				to_sfixed(0.5343,1,L_SIZE),
				to_sfixed(0.5346,1,L_SIZE),
				to_sfixed(0.5349,1,L_SIZE),
				to_sfixed(0.5351,1,L_SIZE),
				to_sfixed(0.5354,1,L_SIZE),
				to_sfixed(0.5356,1,L_SIZE),
				to_sfixed(0.5359,1,L_SIZE),
				to_sfixed(0.5362,1,L_SIZE),
				to_sfixed(0.5364,1,L_SIZE),
				to_sfixed(0.5367,1,L_SIZE),
				to_sfixed(0.5369,1,L_SIZE),
				to_sfixed(0.5372,1,L_SIZE),
				to_sfixed(0.5375,1,L_SIZE),
				to_sfixed(0.5377,1,L_SIZE),
				to_sfixed(0.5380,1,L_SIZE),
				to_sfixed(0.5382,1,L_SIZE),
				to_sfixed(0.5385,1,L_SIZE),
				to_sfixed(0.5388,1,L_SIZE),
				to_sfixed(0.5390,1,L_SIZE),
				to_sfixed(0.5393,1,L_SIZE),
				to_sfixed(0.5395,1,L_SIZE),
				to_sfixed(0.5398,1,L_SIZE),
				to_sfixed(0.5401,1,L_SIZE),
				to_sfixed(0.5403,1,L_SIZE),
				to_sfixed(0.5406,1,L_SIZE),
				to_sfixed(0.5408,1,L_SIZE),
				to_sfixed(0.5411,1,L_SIZE),
				to_sfixed(0.5414,1,L_SIZE),
				to_sfixed(0.5416,1,L_SIZE),
				to_sfixed(0.5419,1,L_SIZE),
				to_sfixed(0.5421,1,L_SIZE),
				to_sfixed(0.5424,1,L_SIZE),
				to_sfixed(0.5427,1,L_SIZE),
				to_sfixed(0.5429,1,L_SIZE),
				to_sfixed(0.5432,1,L_SIZE),
				to_sfixed(0.5434,1,L_SIZE),
				to_sfixed(0.5437,1,L_SIZE),
				to_sfixed(0.5439,1,L_SIZE),
				to_sfixed(0.5442,1,L_SIZE),
				to_sfixed(0.5445,1,L_SIZE),
				to_sfixed(0.5447,1,L_SIZE),
				to_sfixed(0.5450,1,L_SIZE),
				to_sfixed(0.5452,1,L_SIZE),
				to_sfixed(0.5455,1,L_SIZE),
				to_sfixed(0.5457,1,L_SIZE),
				to_sfixed(0.5460,1,L_SIZE),
				to_sfixed(0.5463,1,L_SIZE),
				to_sfixed(0.5465,1,L_SIZE),
				to_sfixed(0.5468,1,L_SIZE),
				to_sfixed(0.5470,1,L_SIZE),
				to_sfixed(0.5473,1,L_SIZE),
				to_sfixed(0.5475,1,L_SIZE),
				to_sfixed(0.5478,1,L_SIZE),
				to_sfixed(0.5481,1,L_SIZE),
				to_sfixed(0.5483,1,L_SIZE),
				to_sfixed(0.5486,1,L_SIZE),
				to_sfixed(0.5488,1,L_SIZE),
				to_sfixed(0.5491,1,L_SIZE),
				to_sfixed(0.5493,1,L_SIZE),
				to_sfixed(0.5496,1,L_SIZE),
				to_sfixed(0.5498,1,L_SIZE),
				to_sfixed(0.5501,1,L_SIZE),
				to_sfixed(0.5504,1,L_SIZE),
				to_sfixed(0.5506,1,L_SIZE),
				to_sfixed(0.5509,1,L_SIZE),
				to_sfixed(0.5511,1,L_SIZE),
				to_sfixed(0.5514,1,L_SIZE),
				to_sfixed(0.5516,1,L_SIZE),
				to_sfixed(0.5519,1,L_SIZE),
				to_sfixed(0.5521,1,L_SIZE),
				to_sfixed(0.5524,1,L_SIZE),
				to_sfixed(0.5527,1,L_SIZE),
				to_sfixed(0.5529,1,L_SIZE),
				to_sfixed(0.5532,1,L_SIZE),
				to_sfixed(0.5534,1,L_SIZE),
				to_sfixed(0.5537,1,L_SIZE),
				to_sfixed(0.5539,1,L_SIZE),
				to_sfixed(0.5542,1,L_SIZE),
				to_sfixed(0.5544,1,L_SIZE),
				to_sfixed(0.5547,1,L_SIZE),
				to_sfixed(0.5549,1,L_SIZE),
				to_sfixed(0.5552,1,L_SIZE),
				to_sfixed(0.5554,1,L_SIZE),
				to_sfixed(0.5557,1,L_SIZE),
				to_sfixed(0.5560,1,L_SIZE),
				to_sfixed(0.5562,1,L_SIZE),
				to_sfixed(0.5565,1,L_SIZE),
				to_sfixed(0.5567,1,L_SIZE),
				to_sfixed(0.5570,1,L_SIZE),
				to_sfixed(0.5572,1,L_SIZE),
				to_sfixed(0.5575,1,L_SIZE),
				to_sfixed(0.5577,1,L_SIZE),
				to_sfixed(0.5580,1,L_SIZE),
				to_sfixed(0.5582,1,L_SIZE),
				to_sfixed(0.5585,1,L_SIZE),
				to_sfixed(0.5587,1,L_SIZE),
				to_sfixed(0.5590,1,L_SIZE),
				to_sfixed(0.5592,1,L_SIZE),
				to_sfixed(0.5595,1,L_SIZE),
				to_sfixed(0.5597,1,L_SIZE),
				to_sfixed(0.5600,1,L_SIZE),
				to_sfixed(0.5602,1,L_SIZE),
				to_sfixed(0.5605,1,L_SIZE),
				to_sfixed(0.5607,1,L_SIZE),
				to_sfixed(0.5610,1,L_SIZE),
				to_sfixed(0.5612,1,L_SIZE),
				to_sfixed(0.5615,1,L_SIZE),
				to_sfixed(0.5617,1,L_SIZE),
				to_sfixed(0.5620,1,L_SIZE),
				to_sfixed(0.5622,1,L_SIZE),
				to_sfixed(0.5625,1,L_SIZE),
				to_sfixed(0.5627,1,L_SIZE),
				to_sfixed(0.5630,1,L_SIZE),
				to_sfixed(0.5632,1,L_SIZE),
				to_sfixed(0.5635,1,L_SIZE),
				to_sfixed(0.5637,1,L_SIZE),
				to_sfixed(0.5640,1,L_SIZE),
				to_sfixed(0.5642,1,L_SIZE),
				to_sfixed(0.5645,1,L_SIZE),
				to_sfixed(0.5647,1,L_SIZE),
				to_sfixed(0.5650,1,L_SIZE),
				to_sfixed(0.5652,1,L_SIZE),
				to_sfixed(0.5655,1,L_SIZE),
				to_sfixed(0.5657,1,L_SIZE),
				to_sfixed(0.5660,1,L_SIZE),
				to_sfixed(0.5662,1,L_SIZE),
				to_sfixed(0.5665,1,L_SIZE),
				to_sfixed(0.5667,1,L_SIZE),
				to_sfixed(0.5670,1,L_SIZE),
				to_sfixed(0.5672,1,L_SIZE),
				to_sfixed(0.5675,1,L_SIZE),
				to_sfixed(0.5677,1,L_SIZE),
				to_sfixed(0.5680,1,L_SIZE),
				to_sfixed(0.5682,1,L_SIZE),
				to_sfixed(0.5685,1,L_SIZE),
				to_sfixed(0.5687,1,L_SIZE),
				to_sfixed(0.5690,1,L_SIZE),
				to_sfixed(0.5692,1,L_SIZE),
				to_sfixed(0.5695,1,L_SIZE),
				to_sfixed(0.5697,1,L_SIZE),
				to_sfixed(0.5700,1,L_SIZE),
				to_sfixed(0.5702,1,L_SIZE),
				to_sfixed(0.5705,1,L_SIZE),
				to_sfixed(0.5707,1,L_SIZE),
				to_sfixed(0.5709,1,L_SIZE),
				to_sfixed(0.5712,1,L_SIZE),
				to_sfixed(0.5714,1,L_SIZE),
				to_sfixed(0.5717,1,L_SIZE),
				to_sfixed(0.5719,1,L_SIZE),
				to_sfixed(0.5722,1,L_SIZE),
				to_sfixed(0.5724,1,L_SIZE),
				to_sfixed(0.5727,1,L_SIZE),
				to_sfixed(0.5729,1,L_SIZE),
				to_sfixed(0.5732,1,L_SIZE),
				to_sfixed(0.5734,1,L_SIZE),
				to_sfixed(0.5737,1,L_SIZE),
				to_sfixed(0.5739,1,L_SIZE),
				to_sfixed(0.5741,1,L_SIZE),
				to_sfixed(0.5744,1,L_SIZE),
				to_sfixed(0.5746,1,L_SIZE),
				to_sfixed(0.5749,1,L_SIZE),
				to_sfixed(0.5751,1,L_SIZE),
				to_sfixed(0.5754,1,L_SIZE),
				to_sfixed(0.5756,1,L_SIZE),
				to_sfixed(0.5759,1,L_SIZE),
				to_sfixed(0.5761,1,L_SIZE),
				to_sfixed(0.5764,1,L_SIZE),
				to_sfixed(0.5766,1,L_SIZE),
				to_sfixed(0.5768,1,L_SIZE),
				to_sfixed(0.5771,1,L_SIZE),
				to_sfixed(0.5773,1,L_SIZE),
				to_sfixed(0.5776,1,L_SIZE),
				to_sfixed(0.5778,1,L_SIZE),
				to_sfixed(0.5781,1,L_SIZE),
				to_sfixed(0.5783,1,L_SIZE),
				to_sfixed(0.5785,1,L_SIZE),
				to_sfixed(0.5788,1,L_SIZE),
				to_sfixed(0.5790,1,L_SIZE),
				to_sfixed(0.5793,1,L_SIZE),
				to_sfixed(0.5795,1,L_SIZE),
				to_sfixed(0.5798,1,L_SIZE),
				to_sfixed(0.5800,1,L_SIZE),
				to_sfixed(0.5803,1,L_SIZE),
				to_sfixed(0.5805,1,L_SIZE),
				to_sfixed(0.5807,1,L_SIZE),
				to_sfixed(0.5810,1,L_SIZE),
				to_sfixed(0.5812,1,L_SIZE),
				to_sfixed(0.5815,1,L_SIZE),
				to_sfixed(0.5817,1,L_SIZE),
				to_sfixed(0.5819,1,L_SIZE),
				to_sfixed(0.5822,1,L_SIZE),
				to_sfixed(0.5824,1,L_SIZE),
				to_sfixed(0.5827,1,L_SIZE),
				to_sfixed(0.5829,1,L_SIZE),
				to_sfixed(0.5832,1,L_SIZE),
				to_sfixed(0.5834,1,L_SIZE),
				to_sfixed(0.5836,1,L_SIZE),
				to_sfixed(0.5839,1,L_SIZE),
				to_sfixed(0.5841,1,L_SIZE),
				to_sfixed(0.5844,1,L_SIZE),
				to_sfixed(0.5846,1,L_SIZE),
				to_sfixed(0.5848,1,L_SIZE),
				to_sfixed(0.5851,1,L_SIZE),
				to_sfixed(0.5853,1,L_SIZE),
				to_sfixed(0.5856,1,L_SIZE),
				to_sfixed(0.5858,1,L_SIZE),
				to_sfixed(0.5861,1,L_SIZE),
				to_sfixed(0.5863,1,L_SIZE),
				to_sfixed(0.5865,1,L_SIZE),
				to_sfixed(0.5868,1,L_SIZE),
				to_sfixed(0.5870,1,L_SIZE),
				to_sfixed(0.5873,1,L_SIZE),
				to_sfixed(0.5875,1,L_SIZE),
				to_sfixed(0.5877,1,L_SIZE),
				to_sfixed(0.5880,1,L_SIZE),
				to_sfixed(0.5882,1,L_SIZE),
				to_sfixed(0.5885,1,L_SIZE),
				to_sfixed(0.5887,1,L_SIZE),
				to_sfixed(0.5889,1,L_SIZE),
				to_sfixed(0.5892,1,L_SIZE),
				to_sfixed(0.5894,1,L_SIZE),
				to_sfixed(0.5896,1,L_SIZE),
				to_sfixed(0.5899,1,L_SIZE),
				to_sfixed(0.5901,1,L_SIZE),
				to_sfixed(0.5904,1,L_SIZE),
				to_sfixed(0.5906,1,L_SIZE),
				to_sfixed(0.5908,1,L_SIZE),
				to_sfixed(0.5911,1,L_SIZE),
				to_sfixed(0.5913,1,L_SIZE),
				to_sfixed(0.5916,1,L_SIZE),
				to_sfixed(0.5918,1,L_SIZE),
				to_sfixed(0.5920,1,L_SIZE),
				to_sfixed(0.5923,1,L_SIZE),
				to_sfixed(0.5925,1,L_SIZE),
				to_sfixed(0.5927,1,L_SIZE),
				to_sfixed(0.5930,1,L_SIZE),
				to_sfixed(0.5932,1,L_SIZE),
				to_sfixed(0.5935,1,L_SIZE),
				to_sfixed(0.5937,1,L_SIZE),
				to_sfixed(0.5939,1,L_SIZE),
				to_sfixed(0.5942,1,L_SIZE),
				to_sfixed(0.5944,1,L_SIZE),
				to_sfixed(0.5946,1,L_SIZE),
				to_sfixed(0.5949,1,L_SIZE),
				to_sfixed(0.5951,1,L_SIZE),
				to_sfixed(0.5954,1,L_SIZE),
				to_sfixed(0.5956,1,L_SIZE),
				to_sfixed(0.5958,1,L_SIZE),
				to_sfixed(0.5961,1,L_SIZE),
				to_sfixed(0.5963,1,L_SIZE),
				to_sfixed(0.5965,1,L_SIZE),
				to_sfixed(0.5968,1,L_SIZE),
				to_sfixed(0.5970,1,L_SIZE),
				to_sfixed(0.5972,1,L_SIZE),
				to_sfixed(0.5975,1,L_SIZE),
				to_sfixed(0.5977,1,L_SIZE),
				to_sfixed(0.5979,1,L_SIZE),
				to_sfixed(0.5982,1,L_SIZE),
				to_sfixed(0.5984,1,L_SIZE),
				to_sfixed(0.5986,1,L_SIZE),
				to_sfixed(0.5989,1,L_SIZE),
				to_sfixed(0.5991,1,L_SIZE),
				to_sfixed(0.5994,1,L_SIZE),
				to_sfixed(0.5996,1,L_SIZE),
				to_sfixed(0.5998,1,L_SIZE),
				to_sfixed(0.6001,1,L_SIZE),
				to_sfixed(0.6003,1,L_SIZE),
				to_sfixed(0.6005,1,L_SIZE),
				to_sfixed(0.6008,1,L_SIZE),
				to_sfixed(0.6010,1,L_SIZE),
				to_sfixed(0.6012,1,L_SIZE),
				to_sfixed(0.6015,1,L_SIZE),
				to_sfixed(0.6017,1,L_SIZE),
				to_sfixed(0.6019,1,L_SIZE),
				to_sfixed(0.6022,1,L_SIZE),
				to_sfixed(0.6024,1,L_SIZE),
				to_sfixed(0.6026,1,L_SIZE),
				to_sfixed(0.6029,1,L_SIZE),
				to_sfixed(0.6031,1,L_SIZE),
				to_sfixed(0.6033,1,L_SIZE),
				to_sfixed(0.6036,1,L_SIZE),
				to_sfixed(0.6038,1,L_SIZE),
				to_sfixed(0.6040,1,L_SIZE),
				to_sfixed(0.6043,1,L_SIZE),
				to_sfixed(0.6045,1,L_SIZE),
				to_sfixed(0.6047,1,L_SIZE),
				to_sfixed(0.6050,1,L_SIZE),
				to_sfixed(0.6052,1,L_SIZE),
				to_sfixed(0.6054,1,L_SIZE),
				to_sfixed(0.6057,1,L_SIZE),
				to_sfixed(0.6059,1,L_SIZE),
				to_sfixed(0.6061,1,L_SIZE),
				to_sfixed(0.6063,1,L_SIZE),
				to_sfixed(0.6066,1,L_SIZE),
				to_sfixed(0.6068,1,L_SIZE),
				to_sfixed(0.6070,1,L_SIZE),
				to_sfixed(0.6073,1,L_SIZE),
				to_sfixed(0.6075,1,L_SIZE),
				to_sfixed(0.6077,1,L_SIZE),
				to_sfixed(0.6080,1,L_SIZE),
				to_sfixed(0.6082,1,L_SIZE),
				to_sfixed(0.6084,1,L_SIZE),
				to_sfixed(0.6087,1,L_SIZE),
				to_sfixed(0.6089,1,L_SIZE),
				to_sfixed(0.6091,1,L_SIZE),
				to_sfixed(0.6093,1,L_SIZE),
				to_sfixed(0.6096,1,L_SIZE),
				to_sfixed(0.6098,1,L_SIZE),
				to_sfixed(0.6100,1,L_SIZE),
				to_sfixed(0.6103,1,L_SIZE),
				to_sfixed(0.6105,1,L_SIZE),
				to_sfixed(0.6107,1,L_SIZE),
				to_sfixed(0.6110,1,L_SIZE),
				to_sfixed(0.6112,1,L_SIZE),
				to_sfixed(0.6114,1,L_SIZE),
				to_sfixed(0.6116,1,L_SIZE),
				to_sfixed(0.6119,1,L_SIZE),
				to_sfixed(0.6121,1,L_SIZE),
				to_sfixed(0.6123,1,L_SIZE),
				to_sfixed(0.6126,1,L_SIZE),
				to_sfixed(0.6128,1,L_SIZE),
				to_sfixed(0.6130,1,L_SIZE),
				to_sfixed(0.6132,1,L_SIZE),
				to_sfixed(0.6135,1,L_SIZE),
				to_sfixed(0.6137,1,L_SIZE),
				to_sfixed(0.6139,1,L_SIZE),
				to_sfixed(0.6142,1,L_SIZE),
				to_sfixed(0.6144,1,L_SIZE),
				to_sfixed(0.6146,1,L_SIZE),
				to_sfixed(0.6148,1,L_SIZE),
				to_sfixed(0.6151,1,L_SIZE),
				to_sfixed(0.6153,1,L_SIZE),
				to_sfixed(0.6155,1,L_SIZE),
				to_sfixed(0.6158,1,L_SIZE),
				to_sfixed(0.6160,1,L_SIZE),
				to_sfixed(0.6162,1,L_SIZE),
				to_sfixed(0.6164,1,L_SIZE),
				to_sfixed(0.6167,1,L_SIZE),
				to_sfixed(0.6169,1,L_SIZE),
				to_sfixed(0.6171,1,L_SIZE),
				to_sfixed(0.6173,1,L_SIZE),
				to_sfixed(0.6176,1,L_SIZE),
				to_sfixed(0.6178,1,L_SIZE),
				to_sfixed(0.6180,1,L_SIZE),
				to_sfixed(0.6183,1,L_SIZE),
				to_sfixed(0.6185,1,L_SIZE),
				to_sfixed(0.6187,1,L_SIZE),
				to_sfixed(0.6189,1,L_SIZE),
				to_sfixed(0.6192,1,L_SIZE),
				to_sfixed(0.6194,1,L_SIZE),
				to_sfixed(0.6196,1,L_SIZE),
				to_sfixed(0.6198,1,L_SIZE),
				to_sfixed(0.6201,1,L_SIZE),
				to_sfixed(0.6203,1,L_SIZE),
				to_sfixed(0.6205,1,L_SIZE),
				to_sfixed(0.6207,1,L_SIZE),
				to_sfixed(0.6210,1,L_SIZE),
				to_sfixed(0.6212,1,L_SIZE),
				to_sfixed(0.6214,1,L_SIZE),
				to_sfixed(0.6216,1,L_SIZE),
				to_sfixed(0.6219,1,L_SIZE),
				to_sfixed(0.6221,1,L_SIZE),
				to_sfixed(0.6223,1,L_SIZE),
				to_sfixed(0.6225,1,L_SIZE),
				to_sfixed(0.6228,1,L_SIZE),
				to_sfixed(0.6230,1,L_SIZE),
				to_sfixed(0.6232,1,L_SIZE),
				to_sfixed(0.6234,1,L_SIZE),
				to_sfixed(0.6237,1,L_SIZE),
				to_sfixed(0.6239,1,L_SIZE),
				to_sfixed(0.6241,1,L_SIZE),
				to_sfixed(0.6243,1,L_SIZE),
				to_sfixed(0.6245,1,L_SIZE),
				to_sfixed(0.6248,1,L_SIZE),
				to_sfixed(0.6250,1,L_SIZE),
				to_sfixed(0.6252,1,L_SIZE),
				to_sfixed(0.6254,1,L_SIZE),
				to_sfixed(0.6257,1,L_SIZE),
				to_sfixed(0.6259,1,L_SIZE),
				to_sfixed(0.6261,1,L_SIZE),
				to_sfixed(0.6263,1,L_SIZE),
				to_sfixed(0.6266,1,L_SIZE),
				to_sfixed(0.6268,1,L_SIZE),
				to_sfixed(0.6270,1,L_SIZE),
				to_sfixed(0.6272,1,L_SIZE),
				to_sfixed(0.6274,1,L_SIZE),
				to_sfixed(0.6277,1,L_SIZE),
				to_sfixed(0.6279,1,L_SIZE),
				to_sfixed(0.6281,1,L_SIZE),
				to_sfixed(0.6283,1,L_SIZE),
				to_sfixed(0.6285,1,L_SIZE),
				to_sfixed(0.6288,1,L_SIZE),
				to_sfixed(0.6290,1,L_SIZE),
				to_sfixed(0.6292,1,L_SIZE),
				to_sfixed(0.6294,1,L_SIZE),
				to_sfixed(0.6297,1,L_SIZE),
				to_sfixed(0.6299,1,L_SIZE),
				to_sfixed(0.6301,1,L_SIZE),
				to_sfixed(0.6303,1,L_SIZE),
				to_sfixed(0.6305,1,L_SIZE),
				to_sfixed(0.6308,1,L_SIZE),
				to_sfixed(0.6310,1,L_SIZE),
				to_sfixed(0.6312,1,L_SIZE),
				to_sfixed(0.6314,1,L_SIZE),
				to_sfixed(0.6316,1,L_SIZE),
				to_sfixed(0.6319,1,L_SIZE),
				to_sfixed(0.6321,1,L_SIZE),
				to_sfixed(0.6323,1,L_SIZE),
				to_sfixed(0.6325,1,L_SIZE),
				to_sfixed(0.6327,1,L_SIZE),
				to_sfixed(0.6330,1,L_SIZE),
				to_sfixed(0.6332,1,L_SIZE),
				to_sfixed(0.6334,1,L_SIZE),
				to_sfixed(0.6336,1,L_SIZE),
				to_sfixed(0.6338,1,L_SIZE),
				to_sfixed(0.6341,1,L_SIZE),
				to_sfixed(0.6343,1,L_SIZE),
				to_sfixed(0.6345,1,L_SIZE),
				to_sfixed(0.6347,1,L_SIZE),
				to_sfixed(0.6349,1,L_SIZE),
				to_sfixed(0.6351,1,L_SIZE),
				to_sfixed(0.6354,1,L_SIZE),
				to_sfixed(0.6356,1,L_SIZE),
				to_sfixed(0.6358,1,L_SIZE),
				to_sfixed(0.6360,1,L_SIZE),
				to_sfixed(0.6362,1,L_SIZE),
				to_sfixed(0.6365,1,L_SIZE),
				to_sfixed(0.6367,1,L_SIZE),
				to_sfixed(0.6369,1,L_SIZE),
				to_sfixed(0.6371,1,L_SIZE),
				to_sfixed(0.6373,1,L_SIZE),
				to_sfixed(0.6375,1,L_SIZE),
				to_sfixed(0.6378,1,L_SIZE),
				to_sfixed(0.6380,1,L_SIZE),
				to_sfixed(0.6382,1,L_SIZE),
				to_sfixed(0.6384,1,L_SIZE),
				to_sfixed(0.6386,1,L_SIZE),
				to_sfixed(0.6388,1,L_SIZE),
				to_sfixed(0.6391,1,L_SIZE),
				to_sfixed(0.6393,1,L_SIZE),
				to_sfixed(0.6395,1,L_SIZE),
				to_sfixed(0.6397,1,L_SIZE),
				to_sfixed(0.6399,1,L_SIZE),
				to_sfixed(0.6401,1,L_SIZE),
				to_sfixed(0.6404,1,L_SIZE),
				to_sfixed(0.6406,1,L_SIZE),
				to_sfixed(0.6408,1,L_SIZE),
				to_sfixed(0.6410,1,L_SIZE),
				to_sfixed(0.6412,1,L_SIZE),
				to_sfixed(0.6414,1,L_SIZE),
				to_sfixed(0.6417,1,L_SIZE),
				to_sfixed(0.6419,1,L_SIZE),
				to_sfixed(0.6421,1,L_SIZE),
				to_sfixed(0.6423,1,L_SIZE),
				to_sfixed(0.6425,1,L_SIZE),
				to_sfixed(0.6427,1,L_SIZE),
				to_sfixed(0.6429,1,L_SIZE),
				to_sfixed(0.6432,1,L_SIZE),
				to_sfixed(0.6434,1,L_SIZE),
				to_sfixed(0.6436,1,L_SIZE),
				to_sfixed(0.6438,1,L_SIZE),
				to_sfixed(0.6440,1,L_SIZE),
				to_sfixed(0.6442,1,L_SIZE),
				to_sfixed(0.6444,1,L_SIZE),
				to_sfixed(0.6447,1,L_SIZE),
				to_sfixed(0.6449,1,L_SIZE),
				to_sfixed(0.6451,1,L_SIZE),
				to_sfixed(0.6453,1,L_SIZE),
				to_sfixed(0.6455,1,L_SIZE),
				to_sfixed(0.6457,1,L_SIZE),
				to_sfixed(0.6459,1,L_SIZE),
				to_sfixed(0.6462,1,L_SIZE),
				to_sfixed(0.6464,1,L_SIZE),
				to_sfixed(0.6466,1,L_SIZE),
				to_sfixed(0.6468,1,L_SIZE),
				to_sfixed(0.6470,1,L_SIZE),
				to_sfixed(0.6472,1,L_SIZE),
				to_sfixed(0.6474,1,L_SIZE),
				to_sfixed(0.6477,1,L_SIZE),
				to_sfixed(0.6479,1,L_SIZE),
				to_sfixed(0.6481,1,L_SIZE),
				to_sfixed(0.6483,1,L_SIZE),
				to_sfixed(0.6485,1,L_SIZE),
				to_sfixed(0.6487,1,L_SIZE),
				to_sfixed(0.6489,1,L_SIZE),
				to_sfixed(0.6491,1,L_SIZE),
				to_sfixed(0.6493,1,L_SIZE),
				to_sfixed(0.6496,1,L_SIZE),
				to_sfixed(0.6498,1,L_SIZE),
				to_sfixed(0.6500,1,L_SIZE),
				to_sfixed(0.6502,1,L_SIZE),
				to_sfixed(0.6504,1,L_SIZE),
				to_sfixed(0.6506,1,L_SIZE),
				to_sfixed(0.6508,1,L_SIZE),
				to_sfixed(0.6510,1,L_SIZE),
				to_sfixed(0.6512,1,L_SIZE),
				to_sfixed(0.6515,1,L_SIZE),
				to_sfixed(0.6517,1,L_SIZE),
				to_sfixed(0.6519,1,L_SIZE),
				to_sfixed(0.6521,1,L_SIZE),
				to_sfixed(0.6523,1,L_SIZE),
				to_sfixed(0.6525,1,L_SIZE),
				to_sfixed(0.6527,1,L_SIZE),
				to_sfixed(0.6529,1,L_SIZE),
				to_sfixed(0.6531,1,L_SIZE),
				to_sfixed(0.6534,1,L_SIZE),
				to_sfixed(0.6536,1,L_SIZE),
				to_sfixed(0.6538,1,L_SIZE),
				to_sfixed(0.6540,1,L_SIZE),
				to_sfixed(0.6542,1,L_SIZE),
				to_sfixed(0.6544,1,L_SIZE),
				to_sfixed(0.6546,1,L_SIZE),
				to_sfixed(0.6548,1,L_SIZE),
				to_sfixed(0.6550,1,L_SIZE),
				to_sfixed(0.6552,1,L_SIZE),
				to_sfixed(0.6554,1,L_SIZE),
				to_sfixed(0.6557,1,L_SIZE),
				to_sfixed(0.6559,1,L_SIZE),
				to_sfixed(0.6561,1,L_SIZE),
				to_sfixed(0.6563,1,L_SIZE),
				to_sfixed(0.6565,1,L_SIZE),
				to_sfixed(0.6567,1,L_SIZE),
				to_sfixed(0.6569,1,L_SIZE),
				to_sfixed(0.6571,1,L_SIZE),
				to_sfixed(0.6573,1,L_SIZE),
				to_sfixed(0.6575,1,L_SIZE),
				to_sfixed(0.6577,1,L_SIZE),
				to_sfixed(0.6579,1,L_SIZE),
				to_sfixed(0.6582,1,L_SIZE),
				to_sfixed(0.6584,1,L_SIZE),
				to_sfixed(0.6586,1,L_SIZE),
				to_sfixed(0.6588,1,L_SIZE),
				to_sfixed(0.6590,1,L_SIZE),
				to_sfixed(0.6592,1,L_SIZE),
				to_sfixed(0.6594,1,L_SIZE),
				to_sfixed(0.6596,1,L_SIZE),
				to_sfixed(0.6598,1,L_SIZE),
				to_sfixed(0.6600,1,L_SIZE),
				to_sfixed(0.6602,1,L_SIZE),
				to_sfixed(0.6604,1,L_SIZE),
				to_sfixed(0.6606,1,L_SIZE),
				to_sfixed(0.6608,1,L_SIZE),
				to_sfixed(0.6611,1,L_SIZE),
				to_sfixed(0.6613,1,L_SIZE),
				to_sfixed(0.6615,1,L_SIZE),
				to_sfixed(0.6617,1,L_SIZE),
				to_sfixed(0.6619,1,L_SIZE),
				to_sfixed(0.6621,1,L_SIZE),
				to_sfixed(0.6623,1,L_SIZE),
				to_sfixed(0.6625,1,L_SIZE),
				to_sfixed(0.6627,1,L_SIZE),
				to_sfixed(0.6629,1,L_SIZE),
				to_sfixed(0.6631,1,L_SIZE),
				to_sfixed(0.6633,1,L_SIZE),
				to_sfixed(0.6635,1,L_SIZE),
				to_sfixed(0.6637,1,L_SIZE),
				to_sfixed(0.6639,1,L_SIZE),
				to_sfixed(0.6641,1,L_SIZE),
				to_sfixed(0.6643,1,L_SIZE),
				to_sfixed(0.6645,1,L_SIZE),
				to_sfixed(0.6647,1,L_SIZE),
				to_sfixed(0.6650,1,L_SIZE),
				to_sfixed(0.6652,1,L_SIZE),
				to_sfixed(0.6654,1,L_SIZE),
				to_sfixed(0.6656,1,L_SIZE),
				to_sfixed(0.6658,1,L_SIZE),
				to_sfixed(0.6660,1,L_SIZE),
				to_sfixed(0.6662,1,L_SIZE),
				to_sfixed(0.6664,1,L_SIZE),
				to_sfixed(0.6666,1,L_SIZE),
				to_sfixed(0.6668,1,L_SIZE),
				to_sfixed(0.6670,1,L_SIZE),
				to_sfixed(0.6672,1,L_SIZE),
				to_sfixed(0.6674,1,L_SIZE),
				to_sfixed(0.6676,1,L_SIZE),
				to_sfixed(0.6678,1,L_SIZE),
				to_sfixed(0.6680,1,L_SIZE),
				to_sfixed(0.6682,1,L_SIZE),
				to_sfixed(0.6684,1,L_SIZE),
				to_sfixed(0.6686,1,L_SIZE),
				to_sfixed(0.6688,1,L_SIZE),
				to_sfixed(0.6690,1,L_SIZE),
				to_sfixed(0.6692,1,L_SIZE),
				to_sfixed(0.6694,1,L_SIZE),
				to_sfixed(0.6696,1,L_SIZE),
				to_sfixed(0.6698,1,L_SIZE),
				to_sfixed(0.6700,1,L_SIZE),
				to_sfixed(0.6702,1,L_SIZE),
				to_sfixed(0.6704,1,L_SIZE),
				to_sfixed(0.6706,1,L_SIZE),
				to_sfixed(0.6708,1,L_SIZE),
				to_sfixed(0.6710,1,L_SIZE),
				to_sfixed(0.6712,1,L_SIZE),
				to_sfixed(0.6714,1,L_SIZE),
				to_sfixed(0.6716,1,L_SIZE),
				to_sfixed(0.6718,1,L_SIZE),
				to_sfixed(0.6720,1,L_SIZE),
				to_sfixed(0.6722,1,L_SIZE),
				to_sfixed(0.6724,1,L_SIZE),
				to_sfixed(0.6726,1,L_SIZE),
				to_sfixed(0.6728,1,L_SIZE),
				to_sfixed(0.6730,1,L_SIZE),
				to_sfixed(0.6732,1,L_SIZE),
				to_sfixed(0.6734,1,L_SIZE),
				to_sfixed(0.6736,1,L_SIZE),
				to_sfixed(0.6738,1,L_SIZE),
				to_sfixed(0.6740,1,L_SIZE),
				to_sfixed(0.6742,1,L_SIZE),
				to_sfixed(0.6744,1,L_SIZE),
				to_sfixed(0.6746,1,L_SIZE),
				to_sfixed(0.6748,1,L_SIZE),
				to_sfixed(0.6750,1,L_SIZE),
				to_sfixed(0.6752,1,L_SIZE),
				to_sfixed(0.6754,1,L_SIZE),
				to_sfixed(0.6756,1,L_SIZE),
				to_sfixed(0.6758,1,L_SIZE),
				to_sfixed(0.6760,1,L_SIZE),
				to_sfixed(0.6762,1,L_SIZE),
				to_sfixed(0.6764,1,L_SIZE),
				to_sfixed(0.6766,1,L_SIZE),
				to_sfixed(0.6768,1,L_SIZE),
				to_sfixed(0.6770,1,L_SIZE),
				to_sfixed(0.6772,1,L_SIZE),
				to_sfixed(0.6774,1,L_SIZE),
				to_sfixed(0.6776,1,L_SIZE),
				to_sfixed(0.6778,1,L_SIZE),
				to_sfixed(0.6780,1,L_SIZE),
				to_sfixed(0.6782,1,L_SIZE),
				to_sfixed(0.6784,1,L_SIZE),
				to_sfixed(0.6786,1,L_SIZE),
				to_sfixed(0.6788,1,L_SIZE),
				to_sfixed(0.6790,1,L_SIZE),
				to_sfixed(0.6792,1,L_SIZE),
				to_sfixed(0.6794,1,L_SIZE),
				to_sfixed(0.6796,1,L_SIZE),
				to_sfixed(0.6798,1,L_SIZE),
				to_sfixed(0.6800,1,L_SIZE),
				to_sfixed(0.6802,1,L_SIZE),
				to_sfixed(0.6804,1,L_SIZE),
				to_sfixed(0.6806,1,L_SIZE),
				to_sfixed(0.6808,1,L_SIZE),
				to_sfixed(0.6810,1,L_SIZE),
				to_sfixed(0.6812,1,L_SIZE),
				to_sfixed(0.6814,1,L_SIZE),
				to_sfixed(0.6816,1,L_SIZE),
				to_sfixed(0.6818,1,L_SIZE),
				to_sfixed(0.6820,1,L_SIZE),
				to_sfixed(0.6822,1,L_SIZE),
				to_sfixed(0.6823,1,L_SIZE),
				to_sfixed(0.6825,1,L_SIZE),
				to_sfixed(0.6827,1,L_SIZE),
				to_sfixed(0.6829,1,L_SIZE),
				to_sfixed(0.6831,1,L_SIZE),
				to_sfixed(0.6833,1,L_SIZE),
				to_sfixed(0.6835,1,L_SIZE),
				to_sfixed(0.6837,1,L_SIZE),
				to_sfixed(0.6839,1,L_SIZE),
				to_sfixed(0.6841,1,L_SIZE),
				to_sfixed(0.6843,1,L_SIZE),
				to_sfixed(0.6845,1,L_SIZE),
				to_sfixed(0.6847,1,L_SIZE),
				to_sfixed(0.6849,1,L_SIZE),
				to_sfixed(0.6851,1,L_SIZE),
				to_sfixed(0.6853,1,L_SIZE),
				to_sfixed(0.6855,1,L_SIZE),
				to_sfixed(0.6857,1,L_SIZE),
				to_sfixed(0.6859,1,L_SIZE),
				to_sfixed(0.6860,1,L_SIZE),
				to_sfixed(0.6862,1,L_SIZE),
				to_sfixed(0.6864,1,L_SIZE),
				to_sfixed(0.6866,1,L_SIZE),
				to_sfixed(0.6868,1,L_SIZE),
				to_sfixed(0.6870,1,L_SIZE),
				to_sfixed(0.6872,1,L_SIZE),
				to_sfixed(0.6874,1,L_SIZE),
				to_sfixed(0.6876,1,L_SIZE),
				to_sfixed(0.6878,1,L_SIZE),
				to_sfixed(0.6880,1,L_SIZE),
				to_sfixed(0.6882,1,L_SIZE),
				to_sfixed(0.6884,1,L_SIZE),
				to_sfixed(0.6886,1,L_SIZE),
				to_sfixed(0.6888,1,L_SIZE),
				to_sfixed(0.6889,1,L_SIZE),
				to_sfixed(0.6891,1,L_SIZE),
				to_sfixed(0.6893,1,L_SIZE),
				to_sfixed(0.6895,1,L_SIZE),
				to_sfixed(0.6897,1,L_SIZE),
				to_sfixed(0.6899,1,L_SIZE),
				to_sfixed(0.6901,1,L_SIZE),
				to_sfixed(0.6903,1,L_SIZE),
				to_sfixed(0.6905,1,L_SIZE),
				to_sfixed(0.6907,1,L_SIZE),
				to_sfixed(0.6909,1,L_SIZE),
				to_sfixed(0.6911,1,L_SIZE),
				to_sfixed(0.6912,1,L_SIZE),
				to_sfixed(0.6914,1,L_SIZE),
				to_sfixed(0.6916,1,L_SIZE),
				to_sfixed(0.6918,1,L_SIZE),
				to_sfixed(0.6920,1,L_SIZE),
				to_sfixed(0.6922,1,L_SIZE),
				to_sfixed(0.6924,1,L_SIZE),
				to_sfixed(0.6926,1,L_SIZE),
				to_sfixed(0.6928,1,L_SIZE),
				to_sfixed(0.6930,1,L_SIZE),
				to_sfixed(0.6932,1,L_SIZE),
				to_sfixed(0.6933,1,L_SIZE),
				to_sfixed(0.6935,1,L_SIZE),
				to_sfixed(0.6937,1,L_SIZE),
				to_sfixed(0.6939,1,L_SIZE),
				to_sfixed(0.6941,1,L_SIZE),
				to_sfixed(0.6943,1,L_SIZE),
				to_sfixed(0.6945,1,L_SIZE),
				to_sfixed(0.6947,1,L_SIZE),
				to_sfixed(0.6949,1,L_SIZE),
				to_sfixed(0.6951,1,L_SIZE),
				to_sfixed(0.6952,1,L_SIZE),
				to_sfixed(0.6954,1,L_SIZE),
				to_sfixed(0.6956,1,L_SIZE),
				to_sfixed(0.6958,1,L_SIZE),
				to_sfixed(0.6960,1,L_SIZE),
				to_sfixed(0.6962,1,L_SIZE),
				to_sfixed(0.6964,1,L_SIZE),
				to_sfixed(0.6966,1,L_SIZE),
				to_sfixed(0.6968,1,L_SIZE),
				to_sfixed(0.6969,1,L_SIZE),
				to_sfixed(0.6971,1,L_SIZE),
				to_sfixed(0.6973,1,L_SIZE),
				to_sfixed(0.6975,1,L_SIZE),
				to_sfixed(0.6977,1,L_SIZE),
				to_sfixed(0.6979,1,L_SIZE),
				to_sfixed(0.6981,1,L_SIZE),
				to_sfixed(0.6983,1,L_SIZE),
				to_sfixed(0.6984,1,L_SIZE),
				to_sfixed(0.6986,1,L_SIZE),
				to_sfixed(0.6988,1,L_SIZE),
				to_sfixed(0.6990,1,L_SIZE),
				to_sfixed(0.6992,1,L_SIZE),
				to_sfixed(0.6994,1,L_SIZE),
				to_sfixed(0.6996,1,L_SIZE),
				to_sfixed(0.6998,1,L_SIZE),
				to_sfixed(0.6999,1,L_SIZE),
				to_sfixed(0.7001,1,L_SIZE),
				to_sfixed(0.7003,1,L_SIZE),
				to_sfixed(0.7005,1,L_SIZE),
				to_sfixed(0.7007,1,L_SIZE),
				to_sfixed(0.7009,1,L_SIZE),
				to_sfixed(0.7011,1,L_SIZE),
				to_sfixed(0.7012,1,L_SIZE),
				to_sfixed(0.7014,1,L_SIZE),
				to_sfixed(0.7016,1,L_SIZE),
				to_sfixed(0.7018,1,L_SIZE),
				to_sfixed(0.7020,1,L_SIZE),
				to_sfixed(0.7022,1,L_SIZE),
				to_sfixed(0.7024,1,L_SIZE),
				to_sfixed(0.7025,1,L_SIZE),
				to_sfixed(0.7027,1,L_SIZE),
				to_sfixed(0.7029,1,L_SIZE),
				to_sfixed(0.7031,1,L_SIZE),
				to_sfixed(0.7033,1,L_SIZE),
				to_sfixed(0.7035,1,L_SIZE),
				to_sfixed(0.7037,1,L_SIZE),
				to_sfixed(0.7038,1,L_SIZE),
				to_sfixed(0.7040,1,L_SIZE),
				to_sfixed(0.7042,1,L_SIZE),
				to_sfixed(0.7044,1,L_SIZE),
				to_sfixed(0.7046,1,L_SIZE),
				to_sfixed(0.7048,1,L_SIZE),
				to_sfixed(0.7050,1,L_SIZE),
				to_sfixed(0.7051,1,L_SIZE),
				to_sfixed(0.7053,1,L_SIZE),
				to_sfixed(0.7055,1,L_SIZE),
				to_sfixed(0.7057,1,L_SIZE),
				to_sfixed(0.7059,1,L_SIZE),
				to_sfixed(0.7061,1,L_SIZE),
				to_sfixed(0.7062,1,L_SIZE),
				to_sfixed(0.7064,1,L_SIZE),
				to_sfixed(0.7066,1,L_SIZE),
				to_sfixed(0.7068,1,L_SIZE),
				to_sfixed(0.7070,1,L_SIZE),
				to_sfixed(0.7072,1,L_SIZE),
				to_sfixed(0.7073,1,L_SIZE),
				to_sfixed(0.7075,1,L_SIZE),
				to_sfixed(0.7077,1,L_SIZE),
				to_sfixed(0.7079,1,L_SIZE),
				to_sfixed(0.7081,1,L_SIZE),
				to_sfixed(0.7083,1,L_SIZE),
				to_sfixed(0.7084,1,L_SIZE),
				to_sfixed(0.7086,1,L_SIZE),
				to_sfixed(0.7088,1,L_SIZE),
				to_sfixed(0.7090,1,L_SIZE),
				to_sfixed(0.7092,1,L_SIZE),
				to_sfixed(0.7093,1,L_SIZE),
				to_sfixed(0.7095,1,L_SIZE),
				to_sfixed(0.7097,1,L_SIZE),
				to_sfixed(0.7099,1,L_SIZE),
				to_sfixed(0.7101,1,L_SIZE),
				to_sfixed(0.7103,1,L_SIZE),
				to_sfixed(0.7104,1,L_SIZE),
				to_sfixed(0.7106,1,L_SIZE),
				to_sfixed(0.7108,1,L_SIZE),
				to_sfixed(0.7110,1,L_SIZE),
				to_sfixed(0.7112,1,L_SIZE),
				to_sfixed(0.7113,1,L_SIZE),
				to_sfixed(0.7115,1,L_SIZE),
				to_sfixed(0.7117,1,L_SIZE),
				to_sfixed(0.7119,1,L_SIZE),
				to_sfixed(0.7121,1,L_SIZE),
				to_sfixed(0.7122,1,L_SIZE),
				to_sfixed(0.7124,1,L_SIZE),
				to_sfixed(0.7126,1,L_SIZE),
				to_sfixed(0.7128,1,L_SIZE),
				to_sfixed(0.7130,1,L_SIZE),
				to_sfixed(0.7131,1,L_SIZE),
				to_sfixed(0.7133,1,L_SIZE),
				to_sfixed(0.7135,1,L_SIZE),
				to_sfixed(0.7137,1,L_SIZE),
				to_sfixed(0.7139,1,L_SIZE),
				to_sfixed(0.7140,1,L_SIZE),
				to_sfixed(0.7142,1,L_SIZE),
				to_sfixed(0.7144,1,L_SIZE),
				to_sfixed(0.7146,1,L_SIZE),
				to_sfixed(0.7148,1,L_SIZE),
				to_sfixed(0.7149,1,L_SIZE),
				to_sfixed(0.7151,1,L_SIZE),
				to_sfixed(0.7153,1,L_SIZE),
				to_sfixed(0.7155,1,L_SIZE),
				to_sfixed(0.7157,1,L_SIZE),
				to_sfixed(0.7158,1,L_SIZE),
				to_sfixed(0.7160,1,L_SIZE),
				to_sfixed(0.7162,1,L_SIZE),
				to_sfixed(0.7164,1,L_SIZE),
				to_sfixed(0.7165,1,L_SIZE),
				to_sfixed(0.7167,1,L_SIZE),
				to_sfixed(0.7169,1,L_SIZE),
				to_sfixed(0.7171,1,L_SIZE),
				to_sfixed(0.7173,1,L_SIZE),
				to_sfixed(0.7174,1,L_SIZE),
				to_sfixed(0.7176,1,L_SIZE),
				to_sfixed(0.7178,1,L_SIZE),
				to_sfixed(0.7180,1,L_SIZE),
				to_sfixed(0.7181,1,L_SIZE),
				to_sfixed(0.7183,1,L_SIZE),
				to_sfixed(0.7185,1,L_SIZE),
				to_sfixed(0.7187,1,L_SIZE),
				to_sfixed(0.7189,1,L_SIZE),
				to_sfixed(0.7190,1,L_SIZE),
				to_sfixed(0.7192,1,L_SIZE),
				to_sfixed(0.7194,1,L_SIZE),
				to_sfixed(0.7196,1,L_SIZE),
				to_sfixed(0.7197,1,L_SIZE),
				to_sfixed(0.7199,1,L_SIZE),
				to_sfixed(0.7201,1,L_SIZE),
				to_sfixed(0.7203,1,L_SIZE),
				to_sfixed(0.7204,1,L_SIZE),
				to_sfixed(0.7206,1,L_SIZE),
				to_sfixed(0.7208,1,L_SIZE),
				to_sfixed(0.7210,1,L_SIZE),
				to_sfixed(0.7211,1,L_SIZE),
				to_sfixed(0.7213,1,L_SIZE),
				to_sfixed(0.7215,1,L_SIZE),
				to_sfixed(0.7217,1,L_SIZE),
				to_sfixed(0.7219,1,L_SIZE),
				to_sfixed(0.7220,1,L_SIZE),
				to_sfixed(0.7222,1,L_SIZE),
				to_sfixed(0.7224,1,L_SIZE),
				to_sfixed(0.7226,1,L_SIZE),
				to_sfixed(0.7227,1,L_SIZE),
				to_sfixed(0.7229,1,L_SIZE),
				to_sfixed(0.7231,1,L_SIZE),
				to_sfixed(0.7233,1,L_SIZE),
				to_sfixed(0.7234,1,L_SIZE),
				to_sfixed(0.7236,1,L_SIZE),
				to_sfixed(0.7238,1,L_SIZE),
				to_sfixed(0.7239,1,L_SIZE),
				to_sfixed(0.7241,1,L_SIZE),
				to_sfixed(0.7243,1,L_SIZE),
				to_sfixed(0.7245,1,L_SIZE),
				to_sfixed(0.7246,1,L_SIZE),
				to_sfixed(0.7248,1,L_SIZE),
				to_sfixed(0.7250,1,L_SIZE),
				to_sfixed(0.7252,1,L_SIZE),
				to_sfixed(0.7253,1,L_SIZE),
				to_sfixed(0.7255,1,L_SIZE),
				to_sfixed(0.7257,1,L_SIZE),
				to_sfixed(0.7259,1,L_SIZE),
				to_sfixed(0.7260,1,L_SIZE),
				to_sfixed(0.7262,1,L_SIZE),
				to_sfixed(0.7264,1,L_SIZE),
				to_sfixed(0.7266,1,L_SIZE),
				to_sfixed(0.7267,1,L_SIZE),
				to_sfixed(0.7269,1,L_SIZE),
				to_sfixed(0.7271,1,L_SIZE),
				to_sfixed(0.7272,1,L_SIZE),
				to_sfixed(0.7274,1,L_SIZE),
				to_sfixed(0.7276,1,L_SIZE),
				to_sfixed(0.7278,1,L_SIZE),
				to_sfixed(0.7279,1,L_SIZE),
				to_sfixed(0.7281,1,L_SIZE),
				to_sfixed(0.7283,1,L_SIZE),
				to_sfixed(0.7284,1,L_SIZE),
				to_sfixed(0.7286,1,L_SIZE),
				to_sfixed(0.7288,1,L_SIZE),
				to_sfixed(0.7290,1,L_SIZE),
				to_sfixed(0.7291,1,L_SIZE),
				to_sfixed(0.7293,1,L_SIZE),
				to_sfixed(0.7295,1,L_SIZE),
				to_sfixed(0.7297,1,L_SIZE),
				to_sfixed(0.7298,1,L_SIZE),
				to_sfixed(0.7300,1,L_SIZE),
				to_sfixed(0.7302,1,L_SIZE),
				to_sfixed(0.7303,1,L_SIZE),
				to_sfixed(0.7305,1,L_SIZE),
				to_sfixed(0.7307,1,L_SIZE),
				to_sfixed(0.7308,1,L_SIZE),
				to_sfixed(0.7310,1,L_SIZE),
				to_sfixed(0.7312,1,L_SIZE),
				to_sfixed(0.7314,1,L_SIZE),
				to_sfixed(0.7315,1,L_SIZE),
				to_sfixed(0.7317,1,L_SIZE),
				to_sfixed(0.7319,1,L_SIZE),
				to_sfixed(0.7320,1,L_SIZE),
				to_sfixed(0.7322,1,L_SIZE),
				to_sfixed(0.7324,1,L_SIZE),
				to_sfixed(0.7325,1,L_SIZE),
				to_sfixed(0.7327,1,L_SIZE),
				to_sfixed(0.7329,1,L_SIZE),
				to_sfixed(0.7331,1,L_SIZE),
				to_sfixed(0.7332,1,L_SIZE),
				to_sfixed(0.7334,1,L_SIZE),
				to_sfixed(0.7336,1,L_SIZE),
				to_sfixed(0.7337,1,L_SIZE),
				to_sfixed(0.7339,1,L_SIZE),
				to_sfixed(0.7341,1,L_SIZE),
				to_sfixed(0.7342,1,L_SIZE),
				to_sfixed(0.7344,1,L_SIZE),
				to_sfixed(0.7346,1,L_SIZE),
				to_sfixed(0.7347,1,L_SIZE),
				to_sfixed(0.7349,1,L_SIZE),
				to_sfixed(0.7351,1,L_SIZE),
				to_sfixed(0.7353,1,L_SIZE),
				to_sfixed(0.7354,1,L_SIZE),
				to_sfixed(0.7356,1,L_SIZE),
				to_sfixed(0.7358,1,L_SIZE),
				to_sfixed(0.7359,1,L_SIZE),
				to_sfixed(0.7361,1,L_SIZE),
				to_sfixed(0.7363,1,L_SIZE),
				to_sfixed(0.7364,1,L_SIZE),
				to_sfixed(0.7366,1,L_SIZE),
				to_sfixed(0.7368,1,L_SIZE),
				to_sfixed(0.7369,1,L_SIZE),
				to_sfixed(0.7371,1,L_SIZE),
				to_sfixed(0.7373,1,L_SIZE),
				to_sfixed(0.7374,1,L_SIZE),
				to_sfixed(0.7376,1,L_SIZE),
				to_sfixed(0.7378,1,L_SIZE),
				to_sfixed(0.7379,1,L_SIZE),
				to_sfixed(0.7381,1,L_SIZE),
				to_sfixed(0.7383,1,L_SIZE),
				to_sfixed(0.7384,1,L_SIZE),
				to_sfixed(0.7386,1,L_SIZE),
				to_sfixed(0.7388,1,L_SIZE),
				to_sfixed(0.7389,1,L_SIZE),
				to_sfixed(0.7391,1,L_SIZE),
				to_sfixed(0.7393,1,L_SIZE),
				to_sfixed(0.7394,1,L_SIZE),
				to_sfixed(0.7396,1,L_SIZE),
				to_sfixed(0.7398,1,L_SIZE),
				to_sfixed(0.7399,1,L_SIZE),
				to_sfixed(0.7401,1,L_SIZE),
				to_sfixed(0.7403,1,L_SIZE),
				to_sfixed(0.7404,1,L_SIZE),
				to_sfixed(0.7406,1,L_SIZE),
				to_sfixed(0.7408,1,L_SIZE),
				to_sfixed(0.7409,1,L_SIZE),
				to_sfixed(0.7411,1,L_SIZE),
				to_sfixed(0.7412,1,L_SIZE),
				to_sfixed(0.7414,1,L_SIZE),
				to_sfixed(0.7416,1,L_SIZE),
				to_sfixed(0.7417,1,L_SIZE),
				to_sfixed(0.7419,1,L_SIZE),
				to_sfixed(0.7421,1,L_SIZE),
				to_sfixed(0.7422,1,L_SIZE),
				to_sfixed(0.7424,1,L_SIZE),
				to_sfixed(0.7426,1,L_SIZE),
				to_sfixed(0.7427,1,L_SIZE),
				to_sfixed(0.7429,1,L_SIZE),
				to_sfixed(0.7431,1,L_SIZE),
				to_sfixed(0.7432,1,L_SIZE),
				to_sfixed(0.7434,1,L_SIZE),
				to_sfixed(0.7436,1,L_SIZE),
				to_sfixed(0.7437,1,L_SIZE),
				to_sfixed(0.7439,1,L_SIZE),
				to_sfixed(0.7440,1,L_SIZE),
				to_sfixed(0.7442,1,L_SIZE),
				to_sfixed(0.7444,1,L_SIZE),
				to_sfixed(0.7445,1,L_SIZE),
				to_sfixed(0.7447,1,L_SIZE),
				to_sfixed(0.7449,1,L_SIZE),
				to_sfixed(0.7450,1,L_SIZE),
				to_sfixed(0.7452,1,L_SIZE),
				to_sfixed(0.7453,1,L_SIZE),
				to_sfixed(0.7455,1,L_SIZE),
				to_sfixed(0.7457,1,L_SIZE),
				to_sfixed(0.7458,1,L_SIZE),
				to_sfixed(0.7460,1,L_SIZE),
				to_sfixed(0.7462,1,L_SIZE),
				to_sfixed(0.7463,1,L_SIZE),
				to_sfixed(0.7465,1,L_SIZE),
				to_sfixed(0.7466,1,L_SIZE),
				to_sfixed(0.7468,1,L_SIZE),
				to_sfixed(0.7470,1,L_SIZE),
				to_sfixed(0.7471,1,L_SIZE),
				to_sfixed(0.7473,1,L_SIZE),
				to_sfixed(0.7475,1,L_SIZE),
				to_sfixed(0.7476,1,L_SIZE),
				to_sfixed(0.7478,1,L_SIZE),
				to_sfixed(0.7479,1,L_SIZE),
				to_sfixed(0.7481,1,L_SIZE),
				to_sfixed(0.7483,1,L_SIZE),
				to_sfixed(0.7484,1,L_SIZE),
				to_sfixed(0.7486,1,L_SIZE),
				to_sfixed(0.7487,1,L_SIZE),
				to_sfixed(0.7489,1,L_SIZE),
				to_sfixed(0.7491,1,L_SIZE),
				to_sfixed(0.7492,1,L_SIZE),
				to_sfixed(0.7494,1,L_SIZE),
				to_sfixed(0.7495,1,L_SIZE),
				to_sfixed(0.7497,1,L_SIZE),
				to_sfixed(0.7499,1,L_SIZE),
				to_sfixed(0.7500,1,L_SIZE),
				to_sfixed(0.7502,1,L_SIZE),
				to_sfixed(0.7503,1,L_SIZE),
				to_sfixed(0.7505,1,L_SIZE),
				to_sfixed(0.7507,1,L_SIZE),
				to_sfixed(0.7508,1,L_SIZE),
				to_sfixed(0.7510,1,L_SIZE),
				to_sfixed(0.7511,1,L_SIZE),
				to_sfixed(0.7513,1,L_SIZE),
				to_sfixed(0.7515,1,L_SIZE),
				to_sfixed(0.7516,1,L_SIZE),
				to_sfixed(0.7518,1,L_SIZE),
				to_sfixed(0.7519,1,L_SIZE),
				to_sfixed(0.7521,1,L_SIZE),
				to_sfixed(0.7523,1,L_SIZE),
				to_sfixed(0.7524,1,L_SIZE),
				to_sfixed(0.7526,1,L_SIZE),
				to_sfixed(0.7527,1,L_SIZE),
				to_sfixed(0.7529,1,L_SIZE),
				to_sfixed(0.7531,1,L_SIZE),
				to_sfixed(0.7532,1,L_SIZE),
				to_sfixed(0.7534,1,L_SIZE),
				to_sfixed(0.7535,1,L_SIZE),
				to_sfixed(0.7537,1,L_SIZE),
				to_sfixed(0.7538,1,L_SIZE),
				to_sfixed(0.7540,1,L_SIZE),
				to_sfixed(0.7542,1,L_SIZE),
				to_sfixed(0.7543,1,L_SIZE),
				to_sfixed(0.7545,1,L_SIZE),
				to_sfixed(0.7546,1,L_SIZE),
				to_sfixed(0.7548,1,L_SIZE),
				to_sfixed(0.7550,1,L_SIZE),
				to_sfixed(0.7551,1,L_SIZE),
				to_sfixed(0.7553,1,L_SIZE),
				to_sfixed(0.7554,1,L_SIZE),
				to_sfixed(0.7556,1,L_SIZE),
				to_sfixed(0.7557,1,L_SIZE),
				to_sfixed(0.7559,1,L_SIZE),
				to_sfixed(0.7561,1,L_SIZE),
				to_sfixed(0.7562,1,L_SIZE),
				to_sfixed(0.7564,1,L_SIZE),
				to_sfixed(0.7565,1,L_SIZE),
				to_sfixed(0.7567,1,L_SIZE),
				to_sfixed(0.7568,1,L_SIZE),
				to_sfixed(0.7570,1,L_SIZE),
				to_sfixed(0.7571,1,L_SIZE),
				to_sfixed(0.7573,1,L_SIZE),
				to_sfixed(0.7575,1,L_SIZE),
				to_sfixed(0.7576,1,L_SIZE),
				to_sfixed(0.7578,1,L_SIZE),
				to_sfixed(0.7579,1,L_SIZE),
				to_sfixed(0.7581,1,L_SIZE),
				to_sfixed(0.7582,1,L_SIZE),
				to_sfixed(0.7584,1,L_SIZE),
				to_sfixed(0.7586,1,L_SIZE),
				to_sfixed(0.7587,1,L_SIZE),
				to_sfixed(0.7589,1,L_SIZE),
				to_sfixed(0.7590,1,L_SIZE),
				to_sfixed(0.7592,1,L_SIZE),
				to_sfixed(0.7593,1,L_SIZE),
				to_sfixed(0.7595,1,L_SIZE),
				to_sfixed(0.7596,1,L_SIZE),
				to_sfixed(0.7598,1,L_SIZE),
				to_sfixed(0.7599,1,L_SIZE),
				to_sfixed(0.7601,1,L_SIZE),
				to_sfixed(0.7603,1,L_SIZE),
				to_sfixed(0.7604,1,L_SIZE),
				to_sfixed(0.7606,1,L_SIZE),
				to_sfixed(0.7607,1,L_SIZE),
				to_sfixed(0.7609,1,L_SIZE),
				to_sfixed(0.7610,1,L_SIZE),
				to_sfixed(0.7612,1,L_SIZE),
				to_sfixed(0.7613,1,L_SIZE),
				to_sfixed(0.7615,1,L_SIZE),
				to_sfixed(0.7616,1,L_SIZE),
				to_sfixed(0.7618,1,L_SIZE),
				to_sfixed(0.7620,1,L_SIZE),
				to_sfixed(0.7621,1,L_SIZE),
				to_sfixed(0.7623,1,L_SIZE),
				to_sfixed(0.7624,1,L_SIZE),
				to_sfixed(0.7626,1,L_SIZE),
				to_sfixed(0.7627,1,L_SIZE),
				to_sfixed(0.7629,1,L_SIZE),
				to_sfixed(0.7630,1,L_SIZE),
				to_sfixed(0.7632,1,L_SIZE),
				to_sfixed(0.7633,1,L_SIZE),
				to_sfixed(0.7635,1,L_SIZE),
				to_sfixed(0.7636,1,L_SIZE),
				to_sfixed(0.7638,1,L_SIZE),
				to_sfixed(0.7639,1,L_SIZE),
				to_sfixed(0.7641,1,L_SIZE),
				to_sfixed(0.7642,1,L_SIZE),
				to_sfixed(0.7644,1,L_SIZE),
				to_sfixed(0.7646,1,L_SIZE),
				to_sfixed(0.7647,1,L_SIZE),
				to_sfixed(0.7649,1,L_SIZE),
				to_sfixed(0.7650,1,L_SIZE),
				to_sfixed(0.7652,1,L_SIZE),
				to_sfixed(0.7653,1,L_SIZE),
				to_sfixed(0.7655,1,L_SIZE),
				to_sfixed(0.7656,1,L_SIZE),
				to_sfixed(0.7658,1,L_SIZE),
				to_sfixed(0.7659,1,L_SIZE),
				to_sfixed(0.7661,1,L_SIZE),
				to_sfixed(0.7662,1,L_SIZE),
				to_sfixed(0.7664,1,L_SIZE),
				to_sfixed(0.7665,1,L_SIZE),
				to_sfixed(0.7667,1,L_SIZE),
				to_sfixed(0.7668,1,L_SIZE),
				to_sfixed(0.7670,1,L_SIZE),
				to_sfixed(0.7671,1,L_SIZE),
				to_sfixed(0.7673,1,L_SIZE),
				to_sfixed(0.7674,1,L_SIZE),
				to_sfixed(0.7676,1,L_SIZE),
				to_sfixed(0.7677,1,L_SIZE),
				to_sfixed(0.7679,1,L_SIZE),
				to_sfixed(0.7680,1,L_SIZE),
				to_sfixed(0.7682,1,L_SIZE),
				to_sfixed(0.7683,1,L_SIZE),
				to_sfixed(0.7685,1,L_SIZE),
				to_sfixed(0.7686,1,L_SIZE),
				to_sfixed(0.7688,1,L_SIZE),
				to_sfixed(0.7689,1,L_SIZE),
				to_sfixed(0.7691,1,L_SIZE),
				to_sfixed(0.7692,1,L_SIZE),
				to_sfixed(0.7694,1,L_SIZE),
				to_sfixed(0.7695,1,L_SIZE),
				to_sfixed(0.7697,1,L_SIZE),
				to_sfixed(0.7698,1,L_SIZE),
				to_sfixed(0.7700,1,L_SIZE),
				to_sfixed(0.7701,1,L_SIZE),
				to_sfixed(0.7703,1,L_SIZE),
				to_sfixed(0.7704,1,L_SIZE),
				to_sfixed(0.7706,1,L_SIZE),
				to_sfixed(0.7707,1,L_SIZE),
				to_sfixed(0.7709,1,L_SIZE),
				to_sfixed(0.7710,1,L_SIZE),
				to_sfixed(0.7712,1,L_SIZE),
				to_sfixed(0.7713,1,L_SIZE),
				to_sfixed(0.7715,1,L_SIZE),
				to_sfixed(0.7716,1,L_SIZE),
				to_sfixed(0.7718,1,L_SIZE),
				to_sfixed(0.7719,1,L_SIZE),
				to_sfixed(0.7721,1,L_SIZE),
				to_sfixed(0.7722,1,L_SIZE),
				to_sfixed(0.7723,1,L_SIZE),
				to_sfixed(0.7725,1,L_SIZE),
				to_sfixed(0.7726,1,L_SIZE),
				to_sfixed(0.7728,1,L_SIZE),
				to_sfixed(0.7729,1,L_SIZE),
				to_sfixed(0.7731,1,L_SIZE),
				to_sfixed(0.7732,1,L_SIZE),
				to_sfixed(0.7734,1,L_SIZE),
				to_sfixed(0.7735,1,L_SIZE),
				to_sfixed(0.7737,1,L_SIZE),
				to_sfixed(0.7738,1,L_SIZE),
				to_sfixed(0.7740,1,L_SIZE),
				to_sfixed(0.7741,1,L_SIZE),
				to_sfixed(0.7743,1,L_SIZE),
				to_sfixed(0.7744,1,L_SIZE),
				to_sfixed(0.7746,1,L_SIZE),
				to_sfixed(0.7747,1,L_SIZE),
				to_sfixed(0.7748,1,L_SIZE),
				to_sfixed(0.7750,1,L_SIZE),
				to_sfixed(0.7751,1,L_SIZE),
				to_sfixed(0.7753,1,L_SIZE),
				to_sfixed(0.7754,1,L_SIZE),
				to_sfixed(0.7756,1,L_SIZE),
				to_sfixed(0.7757,1,L_SIZE),
				to_sfixed(0.7759,1,L_SIZE),
				to_sfixed(0.7760,1,L_SIZE),
				to_sfixed(0.7762,1,L_SIZE),
				to_sfixed(0.7763,1,L_SIZE),
				to_sfixed(0.7765,1,L_SIZE),
				to_sfixed(0.7766,1,L_SIZE),
				to_sfixed(0.7767,1,L_SIZE),
				to_sfixed(0.7769,1,L_SIZE),
				to_sfixed(0.7770,1,L_SIZE),
				to_sfixed(0.7772,1,L_SIZE),
				to_sfixed(0.7773,1,L_SIZE),
				to_sfixed(0.7775,1,L_SIZE),
				to_sfixed(0.7776,1,L_SIZE),
				to_sfixed(0.7778,1,L_SIZE),
				to_sfixed(0.7779,1,L_SIZE),
				to_sfixed(0.7780,1,L_SIZE),
				to_sfixed(0.7782,1,L_SIZE),
				to_sfixed(0.7783,1,L_SIZE),
				to_sfixed(0.7785,1,L_SIZE),
				to_sfixed(0.7786,1,L_SIZE),
				to_sfixed(0.7788,1,L_SIZE),
				to_sfixed(0.7789,1,L_SIZE),
				to_sfixed(0.7791,1,L_SIZE),
				to_sfixed(0.7792,1,L_SIZE),
				to_sfixed(0.7793,1,L_SIZE),
				to_sfixed(0.7795,1,L_SIZE),
				to_sfixed(0.7796,1,L_SIZE),
				to_sfixed(0.7798,1,L_SIZE),
				to_sfixed(0.7799,1,L_SIZE),
				to_sfixed(0.7801,1,L_SIZE),
				to_sfixed(0.7802,1,L_SIZE),
				to_sfixed(0.7803,1,L_SIZE),
				to_sfixed(0.7805,1,L_SIZE),
				to_sfixed(0.7806,1,L_SIZE),
				to_sfixed(0.7808,1,L_SIZE),
				to_sfixed(0.7809,1,L_SIZE),
				to_sfixed(0.7811,1,L_SIZE),
				to_sfixed(0.7812,1,L_SIZE),
				to_sfixed(0.7814,1,L_SIZE),
				to_sfixed(0.7815,1,L_SIZE),
				to_sfixed(0.7816,1,L_SIZE),
				to_sfixed(0.7818,1,L_SIZE),
				to_sfixed(0.7819,1,L_SIZE),
				to_sfixed(0.7821,1,L_SIZE),
				to_sfixed(0.7822,1,L_SIZE),
				to_sfixed(0.7823,1,L_SIZE),
				to_sfixed(0.7825,1,L_SIZE),
				to_sfixed(0.7826,1,L_SIZE),
				to_sfixed(0.7828,1,L_SIZE),
				to_sfixed(0.7829,1,L_SIZE),
				to_sfixed(0.7831,1,L_SIZE),
				to_sfixed(0.7832,1,L_SIZE),
				to_sfixed(0.7833,1,L_SIZE),
				to_sfixed(0.7835,1,L_SIZE),
				to_sfixed(0.7836,1,L_SIZE),
				to_sfixed(0.7838,1,L_SIZE),
				to_sfixed(0.7839,1,L_SIZE),
				to_sfixed(0.7840,1,L_SIZE),
				to_sfixed(0.7842,1,L_SIZE),
				to_sfixed(0.7843,1,L_SIZE),
				to_sfixed(0.7845,1,L_SIZE),
				to_sfixed(0.7846,1,L_SIZE),
				to_sfixed(0.7848,1,L_SIZE),
				to_sfixed(0.7849,1,L_SIZE),
				to_sfixed(0.7850,1,L_SIZE),
				to_sfixed(0.7852,1,L_SIZE),
				to_sfixed(0.7853,1,L_SIZE),
				to_sfixed(0.7855,1,L_SIZE),
				to_sfixed(0.7856,1,L_SIZE),
				to_sfixed(0.7857,1,L_SIZE),
				to_sfixed(0.7859,1,L_SIZE),
				to_sfixed(0.7860,1,L_SIZE),
				to_sfixed(0.7862,1,L_SIZE),
				to_sfixed(0.7863,1,L_SIZE),
				to_sfixed(0.7864,1,L_SIZE),
				to_sfixed(0.7866,1,L_SIZE),
				to_sfixed(0.7867,1,L_SIZE),
				to_sfixed(0.7869,1,L_SIZE),
				to_sfixed(0.7870,1,L_SIZE),
				to_sfixed(0.7871,1,L_SIZE),
				to_sfixed(0.7873,1,L_SIZE),
				to_sfixed(0.7874,1,L_SIZE),
				to_sfixed(0.7875,1,L_SIZE),
				to_sfixed(0.7877,1,L_SIZE),
				to_sfixed(0.7878,1,L_SIZE),
				to_sfixed(0.7880,1,L_SIZE),
				to_sfixed(0.7881,1,L_SIZE),
				to_sfixed(0.7882,1,L_SIZE),
				to_sfixed(0.7884,1,L_SIZE),
				to_sfixed(0.7885,1,L_SIZE),
				to_sfixed(0.7887,1,L_SIZE),
				to_sfixed(0.7888,1,L_SIZE),
				to_sfixed(0.7889,1,L_SIZE),
				to_sfixed(0.7891,1,L_SIZE),
				to_sfixed(0.7892,1,L_SIZE),
				to_sfixed(0.7893,1,L_SIZE),
				to_sfixed(0.7895,1,L_SIZE),
				to_sfixed(0.7896,1,L_SIZE),
				to_sfixed(0.7898,1,L_SIZE),
				to_sfixed(0.7899,1,L_SIZE),
				to_sfixed(0.7900,1,L_SIZE),
				to_sfixed(0.7902,1,L_SIZE),
				to_sfixed(0.7903,1,L_SIZE),
				to_sfixed(0.7905,1,L_SIZE),
				to_sfixed(0.7906,1,L_SIZE),
				to_sfixed(0.7907,1,L_SIZE),
				to_sfixed(0.7909,1,L_SIZE),
				to_sfixed(0.7910,1,L_SIZE),
				to_sfixed(0.7911,1,L_SIZE),
				to_sfixed(0.7913,1,L_SIZE),
				to_sfixed(0.7914,1,L_SIZE),
				to_sfixed(0.7915,1,L_SIZE),
				to_sfixed(0.7917,1,L_SIZE),
				to_sfixed(0.7918,1,L_SIZE),
				to_sfixed(0.7920,1,L_SIZE),
				to_sfixed(0.7921,1,L_SIZE),
				to_sfixed(0.7922,1,L_SIZE),
				to_sfixed(0.7924,1,L_SIZE),
				to_sfixed(0.7925,1,L_SIZE),
				to_sfixed(0.7926,1,L_SIZE),
				to_sfixed(0.7928,1,L_SIZE),
				to_sfixed(0.7929,1,L_SIZE),
				to_sfixed(0.7930,1,L_SIZE),
				to_sfixed(0.7932,1,L_SIZE),
				to_sfixed(0.7933,1,L_SIZE),
				to_sfixed(0.7935,1,L_SIZE),
				to_sfixed(0.7936,1,L_SIZE),
				to_sfixed(0.7937,1,L_SIZE),
				to_sfixed(0.7939,1,L_SIZE),
				to_sfixed(0.7940,1,L_SIZE),
				to_sfixed(0.7941,1,L_SIZE),
				to_sfixed(0.7943,1,L_SIZE),
				to_sfixed(0.7944,1,L_SIZE),
				to_sfixed(0.7945,1,L_SIZE),
				to_sfixed(0.7947,1,L_SIZE),
				to_sfixed(0.7948,1,L_SIZE),
				to_sfixed(0.7949,1,L_SIZE),
				to_sfixed(0.7951,1,L_SIZE),
				to_sfixed(0.7952,1,L_SIZE),
				to_sfixed(0.7953,1,L_SIZE),
				to_sfixed(0.7955,1,L_SIZE),
				to_sfixed(0.7956,1,L_SIZE),
				to_sfixed(0.7957,1,L_SIZE),
				to_sfixed(0.7959,1,L_SIZE),
				to_sfixed(0.7960,1,L_SIZE),
				to_sfixed(0.7962,1,L_SIZE),
				to_sfixed(0.7963,1,L_SIZE),
				to_sfixed(0.7964,1,L_SIZE),
				to_sfixed(0.7966,1,L_SIZE),
				to_sfixed(0.7967,1,L_SIZE),
				to_sfixed(0.7968,1,L_SIZE),
				to_sfixed(0.7970,1,L_SIZE),
				to_sfixed(0.7971,1,L_SIZE),
				to_sfixed(0.7972,1,L_SIZE),
				to_sfixed(0.7974,1,L_SIZE),
				to_sfixed(0.7975,1,L_SIZE),
				to_sfixed(0.7976,1,L_SIZE),
				to_sfixed(0.7978,1,L_SIZE),
				to_sfixed(0.7979,1,L_SIZE),
				to_sfixed(0.7980,1,L_SIZE),
				to_sfixed(0.7982,1,L_SIZE),
				to_sfixed(0.7983,1,L_SIZE),
				to_sfixed(0.7984,1,L_SIZE),
				to_sfixed(0.7986,1,L_SIZE),
				to_sfixed(0.7987,1,L_SIZE),
				to_sfixed(0.7988,1,L_SIZE),
				to_sfixed(0.7990,1,L_SIZE),
				to_sfixed(0.7991,1,L_SIZE),
				to_sfixed(0.7992,1,L_SIZE),
				to_sfixed(0.7993,1,L_SIZE),
				to_sfixed(0.7995,1,L_SIZE),
				to_sfixed(0.7996,1,L_SIZE),
				to_sfixed(0.7997,1,L_SIZE),
				to_sfixed(0.7999,1,L_SIZE),
				to_sfixed(0.8000,1,L_SIZE),
				to_sfixed(0.8001,1,L_SIZE),
				to_sfixed(0.8003,1,L_SIZE),
				to_sfixed(0.8004,1,L_SIZE),
				to_sfixed(0.8005,1,L_SIZE),
				to_sfixed(0.8007,1,L_SIZE),
				to_sfixed(0.8008,1,L_SIZE),
				to_sfixed(0.8009,1,L_SIZE),
				to_sfixed(0.8011,1,L_SIZE),
				to_sfixed(0.8012,1,L_SIZE),
				to_sfixed(0.8013,1,L_SIZE),
				to_sfixed(0.8015,1,L_SIZE),
				to_sfixed(0.8016,1,L_SIZE),
				to_sfixed(0.8017,1,L_SIZE),
				to_sfixed(0.8018,1,L_SIZE),
				to_sfixed(0.8020,1,L_SIZE),
				to_sfixed(0.8021,1,L_SIZE),
				to_sfixed(0.8022,1,L_SIZE),
				to_sfixed(0.8024,1,L_SIZE),
				to_sfixed(0.8025,1,L_SIZE),
				to_sfixed(0.8026,1,L_SIZE),
				to_sfixed(0.8028,1,L_SIZE),
				to_sfixed(0.8029,1,L_SIZE),
				to_sfixed(0.8030,1,L_SIZE),
				to_sfixed(0.8031,1,L_SIZE),
				to_sfixed(0.8033,1,L_SIZE),
				to_sfixed(0.8034,1,L_SIZE),
				to_sfixed(0.8035,1,L_SIZE),
				to_sfixed(0.8037,1,L_SIZE),
				to_sfixed(0.8038,1,L_SIZE),
				to_sfixed(0.8039,1,L_SIZE),
				to_sfixed(0.8041,1,L_SIZE),
				to_sfixed(0.8042,1,L_SIZE),
				to_sfixed(0.8043,1,L_SIZE),
				to_sfixed(0.8044,1,L_SIZE),
				to_sfixed(0.8046,1,L_SIZE),
				to_sfixed(0.8047,1,L_SIZE),
				to_sfixed(0.8048,1,L_SIZE),
				to_sfixed(0.8050,1,L_SIZE),
				to_sfixed(0.8051,1,L_SIZE),
				to_sfixed(0.8052,1,L_SIZE),
				to_sfixed(0.8053,1,L_SIZE),
				to_sfixed(0.8055,1,L_SIZE),
				to_sfixed(0.8056,1,L_SIZE),
				to_sfixed(0.8057,1,L_SIZE),
				to_sfixed(0.8059,1,L_SIZE),
				to_sfixed(0.8060,1,L_SIZE),
				to_sfixed(0.8061,1,L_SIZE),
				to_sfixed(0.8062,1,L_SIZE),
				to_sfixed(0.8064,1,L_SIZE),
				to_sfixed(0.8065,1,L_SIZE),
				to_sfixed(0.8066,1,L_SIZE),
				to_sfixed(0.8068,1,L_SIZE),
				to_sfixed(0.8069,1,L_SIZE),
				to_sfixed(0.8070,1,L_SIZE),
				to_sfixed(0.8071,1,L_SIZE),
				to_sfixed(0.8073,1,L_SIZE),
				to_sfixed(0.8074,1,L_SIZE),
				to_sfixed(0.8075,1,L_SIZE),
				to_sfixed(0.8077,1,L_SIZE),
				to_sfixed(0.8078,1,L_SIZE),
				to_sfixed(0.8079,1,L_SIZE),
				to_sfixed(0.8080,1,L_SIZE),
				to_sfixed(0.8082,1,L_SIZE),
				to_sfixed(0.8083,1,L_SIZE),
				to_sfixed(0.8084,1,L_SIZE),
				to_sfixed(0.8085,1,L_SIZE),
				to_sfixed(0.8087,1,L_SIZE),
				to_sfixed(0.8088,1,L_SIZE),
				to_sfixed(0.8089,1,L_SIZE),
				to_sfixed(0.8090,1,L_SIZE),
				to_sfixed(0.8092,1,L_SIZE),
				to_sfixed(0.8093,1,L_SIZE),
				to_sfixed(0.8094,1,L_SIZE),
				to_sfixed(0.8096,1,L_SIZE),
				to_sfixed(0.8097,1,L_SIZE),
				to_sfixed(0.8098,1,L_SIZE),
				to_sfixed(0.8099,1,L_SIZE),
				to_sfixed(0.8101,1,L_SIZE),
				to_sfixed(0.8102,1,L_SIZE),
				to_sfixed(0.8103,1,L_SIZE),
				to_sfixed(0.8104,1,L_SIZE),
				to_sfixed(0.8106,1,L_SIZE),
				to_sfixed(0.8107,1,L_SIZE),
				to_sfixed(0.8108,1,L_SIZE),
				to_sfixed(0.8109,1,L_SIZE),
				to_sfixed(0.8111,1,L_SIZE),
				to_sfixed(0.8112,1,L_SIZE),
				to_sfixed(0.8113,1,L_SIZE),
				to_sfixed(0.8114,1,L_SIZE),
				to_sfixed(0.8116,1,L_SIZE),
				to_sfixed(0.8117,1,L_SIZE),
				to_sfixed(0.8118,1,L_SIZE),
				to_sfixed(0.8119,1,L_SIZE),
				to_sfixed(0.8121,1,L_SIZE),
				to_sfixed(0.8122,1,L_SIZE),
				to_sfixed(0.8123,1,L_SIZE),
				to_sfixed(0.8124,1,L_SIZE),
				to_sfixed(0.8126,1,L_SIZE),
				to_sfixed(0.8127,1,L_SIZE),
				to_sfixed(0.8128,1,L_SIZE),
				to_sfixed(0.8129,1,L_SIZE),
				to_sfixed(0.8131,1,L_SIZE),
				to_sfixed(0.8132,1,L_SIZE),
				to_sfixed(0.8133,1,L_SIZE),
				to_sfixed(0.8134,1,L_SIZE),
				to_sfixed(0.8136,1,L_SIZE),
				to_sfixed(0.8137,1,L_SIZE),
				to_sfixed(0.8138,1,L_SIZE),
				to_sfixed(0.8139,1,L_SIZE),
				to_sfixed(0.8140,1,L_SIZE),
				to_sfixed(0.8142,1,L_SIZE),
				to_sfixed(0.8143,1,L_SIZE),
				to_sfixed(0.8144,1,L_SIZE),
				to_sfixed(0.8145,1,L_SIZE),
				to_sfixed(0.8147,1,L_SIZE),
				to_sfixed(0.8148,1,L_SIZE),
				to_sfixed(0.8149,1,L_SIZE),
				to_sfixed(0.8150,1,L_SIZE),
				to_sfixed(0.8152,1,L_SIZE),
				to_sfixed(0.8153,1,L_SIZE),
				to_sfixed(0.8154,1,L_SIZE),
				to_sfixed(0.8155,1,L_SIZE),
				to_sfixed(0.8156,1,L_SIZE),
				to_sfixed(0.8158,1,L_SIZE),
				to_sfixed(0.8159,1,L_SIZE),
				to_sfixed(0.8160,1,L_SIZE),
				to_sfixed(0.8161,1,L_SIZE),
				to_sfixed(0.8163,1,L_SIZE),
				to_sfixed(0.8164,1,L_SIZE),
				to_sfixed(0.8165,1,L_SIZE),
				to_sfixed(0.8166,1,L_SIZE),
				to_sfixed(0.8167,1,L_SIZE),
				to_sfixed(0.8169,1,L_SIZE),
				to_sfixed(0.8170,1,L_SIZE),
				to_sfixed(0.8171,1,L_SIZE),
				to_sfixed(0.8172,1,L_SIZE),
				to_sfixed(0.8174,1,L_SIZE),
				to_sfixed(0.8175,1,L_SIZE),
				to_sfixed(0.8176,1,L_SIZE),
				to_sfixed(0.8177,1,L_SIZE),
				to_sfixed(0.8178,1,L_SIZE),
				to_sfixed(0.8180,1,L_SIZE),
				to_sfixed(0.8181,1,L_SIZE),
				to_sfixed(0.8182,1,L_SIZE),
				to_sfixed(0.8183,1,L_SIZE),
				to_sfixed(0.8184,1,L_SIZE),
				to_sfixed(0.8186,1,L_SIZE),
				to_sfixed(0.8187,1,L_SIZE),
				to_sfixed(0.8188,1,L_SIZE),
				to_sfixed(0.8189,1,L_SIZE),
				to_sfixed(0.8191,1,L_SIZE),
				to_sfixed(0.8192,1,L_SIZE),
				to_sfixed(0.8193,1,L_SIZE),
				to_sfixed(0.8194,1,L_SIZE),
				to_sfixed(0.8195,1,L_SIZE),
				to_sfixed(0.8197,1,L_SIZE),
				to_sfixed(0.8198,1,L_SIZE),
				to_sfixed(0.8199,1,L_SIZE),
				to_sfixed(0.8200,1,L_SIZE),
				to_sfixed(0.8201,1,L_SIZE),
				to_sfixed(0.8203,1,L_SIZE),
				to_sfixed(0.8204,1,L_SIZE),
				to_sfixed(0.8205,1,L_SIZE),
				to_sfixed(0.8206,1,L_SIZE),
				to_sfixed(0.8207,1,L_SIZE),
				to_sfixed(0.8209,1,L_SIZE),
				to_sfixed(0.8210,1,L_SIZE),
				to_sfixed(0.8211,1,L_SIZE),
				to_sfixed(0.8212,1,L_SIZE),
				to_sfixed(0.8213,1,L_SIZE),
				to_sfixed(0.8214,1,L_SIZE),
				to_sfixed(0.8216,1,L_SIZE),
				to_sfixed(0.8217,1,L_SIZE),
				to_sfixed(0.8218,1,L_SIZE),
				to_sfixed(0.8219,1,L_SIZE),
				to_sfixed(0.8220,1,L_SIZE),
				to_sfixed(0.8222,1,L_SIZE),
				to_sfixed(0.8223,1,L_SIZE),
				to_sfixed(0.8224,1,L_SIZE),
				to_sfixed(0.8225,1,L_SIZE),
				to_sfixed(0.8226,1,L_SIZE),
				to_sfixed(0.8228,1,L_SIZE),
				to_sfixed(0.8229,1,L_SIZE),
				to_sfixed(0.8230,1,L_SIZE),
				to_sfixed(0.8231,1,L_SIZE),
				to_sfixed(0.8232,1,L_SIZE),
				to_sfixed(0.8233,1,L_SIZE),
				to_sfixed(0.8235,1,L_SIZE),
				to_sfixed(0.8236,1,L_SIZE),
				to_sfixed(0.8237,1,L_SIZE),
				to_sfixed(0.8238,1,L_SIZE),
				to_sfixed(0.8239,1,L_SIZE),
				to_sfixed(0.8241,1,L_SIZE),
				to_sfixed(0.8242,1,L_SIZE),
				to_sfixed(0.8243,1,L_SIZE),
				to_sfixed(0.8244,1,L_SIZE),
				to_sfixed(0.8245,1,L_SIZE),
				to_sfixed(0.8246,1,L_SIZE),
				to_sfixed(0.8248,1,L_SIZE),
				to_sfixed(0.8249,1,L_SIZE),
				to_sfixed(0.8250,1,L_SIZE),
				to_sfixed(0.8251,1,L_SIZE),
				to_sfixed(0.8252,1,L_SIZE),
				to_sfixed(0.8253,1,L_SIZE),
				to_sfixed(0.8255,1,L_SIZE),
				to_sfixed(0.8256,1,L_SIZE),
				to_sfixed(0.8257,1,L_SIZE),
				to_sfixed(0.8258,1,L_SIZE),
				to_sfixed(0.8259,1,L_SIZE),
				to_sfixed(0.8260,1,L_SIZE),
				to_sfixed(0.8262,1,L_SIZE),
				to_sfixed(0.8263,1,L_SIZE),
				to_sfixed(0.8264,1,L_SIZE),
				to_sfixed(0.8265,1,L_SIZE),
				to_sfixed(0.8266,1,L_SIZE),
				to_sfixed(0.8267,1,L_SIZE),
				to_sfixed(0.8269,1,L_SIZE),
				to_sfixed(0.8270,1,L_SIZE),
				to_sfixed(0.8271,1,L_SIZE),
				to_sfixed(0.8272,1,L_SIZE),
				to_sfixed(0.8273,1,L_SIZE),
				to_sfixed(0.8274,1,L_SIZE),
				to_sfixed(0.8275,1,L_SIZE),
				to_sfixed(0.8277,1,L_SIZE),
				to_sfixed(0.8278,1,L_SIZE),
				to_sfixed(0.8279,1,L_SIZE),
				to_sfixed(0.8280,1,L_SIZE),
				to_sfixed(0.8281,1,L_SIZE),
				to_sfixed(0.8282,1,L_SIZE),
				to_sfixed(0.8284,1,L_SIZE),
				to_sfixed(0.8285,1,L_SIZE),
				to_sfixed(0.8286,1,L_SIZE),
				to_sfixed(0.8287,1,L_SIZE),
				to_sfixed(0.8288,1,L_SIZE),
				to_sfixed(0.8289,1,L_SIZE),
				to_sfixed(0.8290,1,L_SIZE),
				to_sfixed(0.8292,1,L_SIZE),
				to_sfixed(0.8293,1,L_SIZE),
				to_sfixed(0.8294,1,L_SIZE),
				to_sfixed(0.8295,1,L_SIZE),
				to_sfixed(0.8296,1,L_SIZE),
				to_sfixed(0.8297,1,L_SIZE),
				to_sfixed(0.8298,1,L_SIZE),
				to_sfixed(0.8300,1,L_SIZE),
				to_sfixed(0.8301,1,L_SIZE),
				to_sfixed(0.8302,1,L_SIZE),
				to_sfixed(0.8303,1,L_SIZE),
				to_sfixed(0.8304,1,L_SIZE),
				to_sfixed(0.8305,1,L_SIZE),
				to_sfixed(0.8306,1,L_SIZE),
				to_sfixed(0.8307,1,L_SIZE),
				to_sfixed(0.8309,1,L_SIZE),
				to_sfixed(0.8310,1,L_SIZE),
				to_sfixed(0.8311,1,L_SIZE),
				to_sfixed(0.8312,1,L_SIZE),
				to_sfixed(0.8313,1,L_SIZE),
				to_sfixed(0.8314,1,L_SIZE),
				to_sfixed(0.8315,1,L_SIZE),
				to_sfixed(0.8317,1,L_SIZE),
				to_sfixed(0.8318,1,L_SIZE),
				to_sfixed(0.8319,1,L_SIZE),
				to_sfixed(0.8320,1,L_SIZE),
				to_sfixed(0.8321,1,L_SIZE),
				to_sfixed(0.8322,1,L_SIZE),
				to_sfixed(0.8323,1,L_SIZE),
				to_sfixed(0.8324,1,L_SIZE),
				to_sfixed(0.8326,1,L_SIZE),
				to_sfixed(0.8327,1,L_SIZE),
				to_sfixed(0.8328,1,L_SIZE),
				to_sfixed(0.8329,1,L_SIZE),
				to_sfixed(0.8330,1,L_SIZE),
				to_sfixed(0.8331,1,L_SIZE),
				to_sfixed(0.8332,1,L_SIZE),
				to_sfixed(0.8333,1,L_SIZE),
				to_sfixed(0.8335,1,L_SIZE),
				to_sfixed(0.8336,1,L_SIZE),
				to_sfixed(0.8337,1,L_SIZE),
				to_sfixed(0.8338,1,L_SIZE),
				to_sfixed(0.8339,1,L_SIZE),
				to_sfixed(0.8340,1,L_SIZE),
				to_sfixed(0.8341,1,L_SIZE),
				to_sfixed(0.8342,1,L_SIZE),
				to_sfixed(0.8343,1,L_SIZE),
				to_sfixed(0.8345,1,L_SIZE),
				to_sfixed(0.8346,1,L_SIZE),
				to_sfixed(0.8347,1,L_SIZE),
				to_sfixed(0.8348,1,L_SIZE),
				to_sfixed(0.8349,1,L_SIZE),
				to_sfixed(0.8350,1,L_SIZE),
				to_sfixed(0.8351,1,L_SIZE),
				to_sfixed(0.8352,1,L_SIZE),
				to_sfixed(0.8353,1,L_SIZE),
				to_sfixed(0.8355,1,L_SIZE),
				to_sfixed(0.8356,1,L_SIZE),
				to_sfixed(0.8357,1,L_SIZE),
				to_sfixed(0.8358,1,L_SIZE),
				to_sfixed(0.8359,1,L_SIZE),
				to_sfixed(0.8360,1,L_SIZE),
				to_sfixed(0.8361,1,L_SIZE),
				to_sfixed(0.8362,1,L_SIZE),
				to_sfixed(0.8363,1,L_SIZE),
				to_sfixed(0.8364,1,L_SIZE),
				to_sfixed(0.8366,1,L_SIZE),
				to_sfixed(0.8367,1,L_SIZE),
				to_sfixed(0.8368,1,L_SIZE),
				to_sfixed(0.8369,1,L_SIZE),
				to_sfixed(0.8370,1,L_SIZE),
				to_sfixed(0.8371,1,L_SIZE),
				to_sfixed(0.8372,1,L_SIZE),
				to_sfixed(0.8373,1,L_SIZE),
				to_sfixed(0.8374,1,L_SIZE),
				to_sfixed(0.8375,1,L_SIZE),
				to_sfixed(0.8377,1,L_SIZE),
				to_sfixed(0.8378,1,L_SIZE),
				to_sfixed(0.8379,1,L_SIZE),
				to_sfixed(0.8380,1,L_SIZE),
				to_sfixed(0.8381,1,L_SIZE),
				to_sfixed(0.8382,1,L_SIZE),
				to_sfixed(0.8383,1,L_SIZE),
				to_sfixed(0.8384,1,L_SIZE),
				to_sfixed(0.8385,1,L_SIZE),
				to_sfixed(0.8386,1,L_SIZE),
				to_sfixed(0.8387,1,L_SIZE),
				to_sfixed(0.8389,1,L_SIZE),
				to_sfixed(0.8390,1,L_SIZE),
				to_sfixed(0.8391,1,L_SIZE),
				to_sfixed(0.8392,1,L_SIZE),
				to_sfixed(0.8393,1,L_SIZE),
				to_sfixed(0.8394,1,L_SIZE),
				to_sfixed(0.8395,1,L_SIZE),
				to_sfixed(0.8396,1,L_SIZE),
				to_sfixed(0.8397,1,L_SIZE),
				to_sfixed(0.8398,1,L_SIZE),
				to_sfixed(0.8399,1,L_SIZE),
				to_sfixed(0.8400,1,L_SIZE),
				to_sfixed(0.8401,1,L_SIZE),
				to_sfixed(0.8403,1,L_SIZE),
				to_sfixed(0.8404,1,L_SIZE),
				to_sfixed(0.8405,1,L_SIZE),
				to_sfixed(0.8406,1,L_SIZE),
				to_sfixed(0.8407,1,L_SIZE),
				to_sfixed(0.8408,1,L_SIZE),
				to_sfixed(0.8409,1,L_SIZE),
				to_sfixed(0.8410,1,L_SIZE),
				to_sfixed(0.8411,1,L_SIZE),
				to_sfixed(0.8412,1,L_SIZE),
				to_sfixed(0.8413,1,L_SIZE),
				to_sfixed(0.8414,1,L_SIZE),
				to_sfixed(0.8415,1,L_SIZE),
				to_sfixed(0.8417,1,L_SIZE),
				to_sfixed(0.8418,1,L_SIZE),
				to_sfixed(0.8419,1,L_SIZE),
				to_sfixed(0.8420,1,L_SIZE),
				to_sfixed(0.8421,1,L_SIZE),
				to_sfixed(0.8422,1,L_SIZE),
				to_sfixed(0.8423,1,L_SIZE),
				to_sfixed(0.8424,1,L_SIZE),
				to_sfixed(0.8425,1,L_SIZE),
				to_sfixed(0.8426,1,L_SIZE),
				to_sfixed(0.8427,1,L_SIZE),
				to_sfixed(0.8428,1,L_SIZE),
				to_sfixed(0.8429,1,L_SIZE),
				to_sfixed(0.8430,1,L_SIZE),
				to_sfixed(0.8431,1,L_SIZE),
				to_sfixed(0.8432,1,L_SIZE),
				to_sfixed(0.8434,1,L_SIZE),
				to_sfixed(0.8435,1,L_SIZE),
				to_sfixed(0.8436,1,L_SIZE),
				to_sfixed(0.8437,1,L_SIZE),
				to_sfixed(0.8438,1,L_SIZE),
				to_sfixed(0.8439,1,L_SIZE),
				to_sfixed(0.8440,1,L_SIZE),
				to_sfixed(0.8441,1,L_SIZE),
				to_sfixed(0.8442,1,L_SIZE),
				to_sfixed(0.8443,1,L_SIZE),
				to_sfixed(0.8444,1,L_SIZE),
				to_sfixed(0.8445,1,L_SIZE),
				to_sfixed(0.8446,1,L_SIZE),
				to_sfixed(0.8447,1,L_SIZE),
				to_sfixed(0.8448,1,L_SIZE),
				to_sfixed(0.8449,1,L_SIZE),
				to_sfixed(0.8450,1,L_SIZE),
				to_sfixed(0.8451,1,L_SIZE),
				to_sfixed(0.8452,1,L_SIZE),
				to_sfixed(0.8453,1,L_SIZE),
				to_sfixed(0.8455,1,L_SIZE),
				to_sfixed(0.8456,1,L_SIZE),
				to_sfixed(0.8457,1,L_SIZE),
				to_sfixed(0.8458,1,L_SIZE),
				to_sfixed(0.8459,1,L_SIZE),
				to_sfixed(0.8460,1,L_SIZE),
				to_sfixed(0.8461,1,L_SIZE),
				to_sfixed(0.8462,1,L_SIZE),
				to_sfixed(0.8463,1,L_SIZE),
				to_sfixed(0.8464,1,L_SIZE),
				to_sfixed(0.8465,1,L_SIZE),
				to_sfixed(0.8466,1,L_SIZE),
				to_sfixed(0.8467,1,L_SIZE),
				to_sfixed(0.8468,1,L_SIZE),
				to_sfixed(0.8469,1,L_SIZE),
				to_sfixed(0.8470,1,L_SIZE),
				to_sfixed(0.8471,1,L_SIZE),
				to_sfixed(0.8472,1,L_SIZE),
				to_sfixed(0.8473,1,L_SIZE),
				to_sfixed(0.8474,1,L_SIZE),
				to_sfixed(0.8475,1,L_SIZE),
				to_sfixed(0.8476,1,L_SIZE),
				to_sfixed(0.8477,1,L_SIZE),
				to_sfixed(0.8478,1,L_SIZE),
				to_sfixed(0.8479,1,L_SIZE),
				to_sfixed(0.8480,1,L_SIZE),
				to_sfixed(0.8481,1,L_SIZE),
				to_sfixed(0.8482,1,L_SIZE),
				to_sfixed(0.8484,1,L_SIZE),
				to_sfixed(0.8485,1,L_SIZE),
				to_sfixed(0.8486,1,L_SIZE),
				to_sfixed(0.8487,1,L_SIZE),
				to_sfixed(0.8488,1,L_SIZE),
				to_sfixed(0.8489,1,L_SIZE),
				to_sfixed(0.8490,1,L_SIZE),
				to_sfixed(0.8491,1,L_SIZE),
				to_sfixed(0.8492,1,L_SIZE),
				to_sfixed(0.8493,1,L_SIZE),
				to_sfixed(0.8494,1,L_SIZE),
				to_sfixed(0.8495,1,L_SIZE),
				to_sfixed(0.8496,1,L_SIZE),
				to_sfixed(0.8497,1,L_SIZE),
				to_sfixed(0.8498,1,L_SIZE),
				to_sfixed(0.8499,1,L_SIZE),
				to_sfixed(0.8500,1,L_SIZE),
				to_sfixed(0.8501,1,L_SIZE),
				to_sfixed(0.8502,1,L_SIZE),
				to_sfixed(0.8503,1,L_SIZE),
				to_sfixed(0.8504,1,L_SIZE),
				to_sfixed(0.8505,1,L_SIZE),
				to_sfixed(0.8506,1,L_SIZE),
				to_sfixed(0.8507,1,L_SIZE),
				to_sfixed(0.8508,1,L_SIZE),
				to_sfixed(0.8509,1,L_SIZE),
				to_sfixed(0.8510,1,L_SIZE),
				to_sfixed(0.8511,1,L_SIZE),
				to_sfixed(0.8512,1,L_SIZE),
				to_sfixed(0.8513,1,L_SIZE),
				to_sfixed(0.8514,1,L_SIZE),
				to_sfixed(0.8515,1,L_SIZE),
				to_sfixed(0.8516,1,L_SIZE),
				to_sfixed(0.8517,1,L_SIZE),
				to_sfixed(0.8518,1,L_SIZE),
				to_sfixed(0.8519,1,L_SIZE),
				to_sfixed(0.8520,1,L_SIZE),
				to_sfixed(0.8521,1,L_SIZE),
				to_sfixed(0.8522,1,L_SIZE),
				to_sfixed(0.8523,1,L_SIZE),
				to_sfixed(0.8524,1,L_SIZE),
				to_sfixed(0.8525,1,L_SIZE),
				to_sfixed(0.8526,1,L_SIZE),
				to_sfixed(0.8527,1,L_SIZE),
				to_sfixed(0.8528,1,L_SIZE),
				to_sfixed(0.8529,1,L_SIZE),
				to_sfixed(0.8530,1,L_SIZE),
				to_sfixed(0.8531,1,L_SIZE),
				to_sfixed(0.8532,1,L_SIZE),
				to_sfixed(0.8533,1,L_SIZE),
				to_sfixed(0.8534,1,L_SIZE),
				to_sfixed(0.8535,1,L_SIZE),
				to_sfixed(0.8536,1,L_SIZE),
				to_sfixed(0.8537,1,L_SIZE),
				to_sfixed(0.8538,1,L_SIZE),
				to_sfixed(0.8539,1,L_SIZE),
				to_sfixed(0.8540,1,L_SIZE),
				to_sfixed(0.8541,1,L_SIZE),
				to_sfixed(0.8542,1,L_SIZE),
				to_sfixed(0.8543,1,L_SIZE),
				to_sfixed(0.8544,1,L_SIZE),
				to_sfixed(0.8545,1,L_SIZE),
				to_sfixed(0.8546,1,L_SIZE),
				to_sfixed(0.8547,1,L_SIZE),
				to_sfixed(0.8548,1,L_SIZE),
				to_sfixed(0.8549,1,L_SIZE),
				to_sfixed(0.8550,1,L_SIZE),
				to_sfixed(0.8551,1,L_SIZE),
				to_sfixed(0.8552,1,L_SIZE),
				to_sfixed(0.8553,1,L_SIZE),
				to_sfixed(0.8554,1,L_SIZE),
				to_sfixed(0.8555,1,L_SIZE),
				to_sfixed(0.8556,1,L_SIZE),
				to_sfixed(0.8557,1,L_SIZE),
				to_sfixed(0.8558,1,L_SIZE),
				to_sfixed(0.8559,1,L_SIZE),
				to_sfixed(0.8560,1,L_SIZE),
				to_sfixed(0.8561,1,L_SIZE),
				to_sfixed(0.8562,1,L_SIZE),
				to_sfixed(0.8563,1,L_SIZE),
				to_sfixed(0.8564,1,L_SIZE),
				to_sfixed(0.8565,1,L_SIZE),
				to_sfixed(0.8566,1,L_SIZE),
				to_sfixed(0.8567,1,L_SIZE),
				to_sfixed(0.8568,1,L_SIZE),
				to_sfixed(0.8569,1,L_SIZE),
				to_sfixed(0.8569,1,L_SIZE),
				to_sfixed(0.8570,1,L_SIZE),
				to_sfixed(0.8571,1,L_SIZE),
				to_sfixed(0.8572,1,L_SIZE),
				to_sfixed(0.8573,1,L_SIZE),
				to_sfixed(0.8574,1,L_SIZE),
				to_sfixed(0.8575,1,L_SIZE),
				to_sfixed(0.8576,1,L_SIZE),
				to_sfixed(0.8577,1,L_SIZE),
				to_sfixed(0.8578,1,L_SIZE),
				to_sfixed(0.8579,1,L_SIZE),
				to_sfixed(0.8580,1,L_SIZE),
				to_sfixed(0.8581,1,L_SIZE),
				to_sfixed(0.8582,1,L_SIZE),
				to_sfixed(0.8583,1,L_SIZE),
				to_sfixed(0.8584,1,L_SIZE),
				to_sfixed(0.8585,1,L_SIZE),
				to_sfixed(0.8586,1,L_SIZE),
				to_sfixed(0.8587,1,L_SIZE),
				to_sfixed(0.8588,1,L_SIZE),
				to_sfixed(0.8589,1,L_SIZE),
				to_sfixed(0.8590,1,L_SIZE),
				to_sfixed(0.8591,1,L_SIZE),
				to_sfixed(0.8592,1,L_SIZE),
				to_sfixed(0.8593,1,L_SIZE),
				to_sfixed(0.8594,1,L_SIZE),
				to_sfixed(0.8595,1,L_SIZE),
				to_sfixed(0.8596,1,L_SIZE),
				to_sfixed(0.8596,1,L_SIZE),
				to_sfixed(0.8597,1,L_SIZE),
				to_sfixed(0.8598,1,L_SIZE),
				to_sfixed(0.8599,1,L_SIZE),
				to_sfixed(0.8600,1,L_SIZE),
				to_sfixed(0.8601,1,L_SIZE),
				to_sfixed(0.8602,1,L_SIZE),
				to_sfixed(0.8603,1,L_SIZE),
				to_sfixed(0.8604,1,L_SIZE),
				to_sfixed(0.8605,1,L_SIZE),
				to_sfixed(0.8606,1,L_SIZE),
				to_sfixed(0.8607,1,L_SIZE),
				to_sfixed(0.8608,1,L_SIZE),
				to_sfixed(0.8609,1,L_SIZE),
				to_sfixed(0.8610,1,L_SIZE),
				to_sfixed(0.8611,1,L_SIZE),
				to_sfixed(0.8612,1,L_SIZE),
				to_sfixed(0.8613,1,L_SIZE),
				to_sfixed(0.8614,1,L_SIZE),
				to_sfixed(0.8615,1,L_SIZE),
				to_sfixed(0.8615,1,L_SIZE),
				to_sfixed(0.8616,1,L_SIZE),
				to_sfixed(0.8617,1,L_SIZE),
				to_sfixed(0.8618,1,L_SIZE),
				to_sfixed(0.8619,1,L_SIZE),
				to_sfixed(0.8620,1,L_SIZE),
				to_sfixed(0.8621,1,L_SIZE),
				to_sfixed(0.8622,1,L_SIZE),
				to_sfixed(0.8623,1,L_SIZE),
				to_sfixed(0.8624,1,L_SIZE),
				to_sfixed(0.8625,1,L_SIZE),
				to_sfixed(0.8626,1,L_SIZE),
				to_sfixed(0.8627,1,L_SIZE),
				to_sfixed(0.8628,1,L_SIZE),
				to_sfixed(0.8629,1,L_SIZE),
				to_sfixed(0.8630,1,L_SIZE),
				to_sfixed(0.8630,1,L_SIZE),
				to_sfixed(0.8631,1,L_SIZE),
				to_sfixed(0.8632,1,L_SIZE),
				to_sfixed(0.8633,1,L_SIZE),
				to_sfixed(0.8634,1,L_SIZE),
				to_sfixed(0.8635,1,L_SIZE),
				to_sfixed(0.8636,1,L_SIZE),
				to_sfixed(0.8637,1,L_SIZE),
				to_sfixed(0.8638,1,L_SIZE),
				to_sfixed(0.8639,1,L_SIZE),
				to_sfixed(0.8640,1,L_SIZE),
				to_sfixed(0.8641,1,L_SIZE),
				to_sfixed(0.8642,1,L_SIZE),
				to_sfixed(0.8643,1,L_SIZE),
				to_sfixed(0.8644,1,L_SIZE),
				to_sfixed(0.8644,1,L_SIZE),
				to_sfixed(0.8645,1,L_SIZE),
				to_sfixed(0.8646,1,L_SIZE),
				to_sfixed(0.8647,1,L_SIZE),
				to_sfixed(0.8648,1,L_SIZE),
				to_sfixed(0.8649,1,L_SIZE),
				to_sfixed(0.8650,1,L_SIZE),
				to_sfixed(0.8651,1,L_SIZE),
				to_sfixed(0.8652,1,L_SIZE),
				to_sfixed(0.8653,1,L_SIZE),
				to_sfixed(0.8654,1,L_SIZE),
				to_sfixed(0.8655,1,L_SIZE),
				to_sfixed(0.8656,1,L_SIZE),
				to_sfixed(0.8656,1,L_SIZE),
				to_sfixed(0.8657,1,L_SIZE),
				to_sfixed(0.8658,1,L_SIZE),
				to_sfixed(0.8659,1,L_SIZE),
				to_sfixed(0.8660,1,L_SIZE),
				to_sfixed(0.8661,1,L_SIZE),
				to_sfixed(0.8662,1,L_SIZE),
				to_sfixed(0.8663,1,L_SIZE),
				to_sfixed(0.8664,1,L_SIZE),
				to_sfixed(0.8665,1,L_SIZE),
				to_sfixed(0.8666,1,L_SIZE),
				to_sfixed(0.8666,1,L_SIZE),
				to_sfixed(0.8667,1,L_SIZE),
				to_sfixed(0.8668,1,L_SIZE),
				to_sfixed(0.8669,1,L_SIZE),
				to_sfixed(0.8670,1,L_SIZE),
				to_sfixed(0.8671,1,L_SIZE),
				to_sfixed(0.8672,1,L_SIZE),
				to_sfixed(0.8673,1,L_SIZE),
				to_sfixed(0.8674,1,L_SIZE),
				to_sfixed(0.8675,1,L_SIZE),
				to_sfixed(0.8676,1,L_SIZE),
				to_sfixed(0.8676,1,L_SIZE),
				to_sfixed(0.8677,1,L_SIZE),
				to_sfixed(0.8678,1,L_SIZE),
				to_sfixed(0.8679,1,L_SIZE),
				to_sfixed(0.8680,1,L_SIZE),
				to_sfixed(0.8681,1,L_SIZE),
				to_sfixed(0.8682,1,L_SIZE),
				to_sfixed(0.8683,1,L_SIZE),
				to_sfixed(0.8684,1,L_SIZE),
				to_sfixed(0.8685,1,L_SIZE),
				to_sfixed(0.8686,1,L_SIZE),
				to_sfixed(0.8686,1,L_SIZE),
				to_sfixed(0.8687,1,L_SIZE),
				to_sfixed(0.8688,1,L_SIZE),
				to_sfixed(0.8689,1,L_SIZE),
				to_sfixed(0.8690,1,L_SIZE),
				to_sfixed(0.8691,1,L_SIZE),
				to_sfixed(0.8692,1,L_SIZE),
				to_sfixed(0.8693,1,L_SIZE),
				to_sfixed(0.8694,1,L_SIZE),
				to_sfixed(0.8694,1,L_SIZE),
				to_sfixed(0.8695,1,L_SIZE),
				to_sfixed(0.8696,1,L_SIZE),
				to_sfixed(0.8697,1,L_SIZE),
				to_sfixed(0.8698,1,L_SIZE),
				to_sfixed(0.8699,1,L_SIZE),
				to_sfixed(0.8700,1,L_SIZE),
				to_sfixed(0.8701,1,L_SIZE),
				to_sfixed(0.8702,1,L_SIZE),
				to_sfixed(0.8702,1,L_SIZE),
				to_sfixed(0.8703,1,L_SIZE),
				to_sfixed(0.8704,1,L_SIZE),
				to_sfixed(0.8705,1,L_SIZE),
				to_sfixed(0.8706,1,L_SIZE),
				to_sfixed(0.8707,1,L_SIZE),
				to_sfixed(0.8708,1,L_SIZE),
				to_sfixed(0.8709,1,L_SIZE),
				to_sfixed(0.8710,1,L_SIZE),
				to_sfixed(0.8710,1,L_SIZE),
				to_sfixed(0.8711,1,L_SIZE),
				to_sfixed(0.8712,1,L_SIZE),
				to_sfixed(0.8713,1,L_SIZE),
				to_sfixed(0.8714,1,L_SIZE),
				to_sfixed(0.8715,1,L_SIZE),
				to_sfixed(0.8716,1,L_SIZE),
				to_sfixed(0.8717,1,L_SIZE),
				to_sfixed(0.8718,1,L_SIZE),
				to_sfixed(0.8718,1,L_SIZE),
				to_sfixed(0.8719,1,L_SIZE),
				to_sfixed(0.8720,1,L_SIZE),
				to_sfixed(0.8721,1,L_SIZE),
				to_sfixed(0.8722,1,L_SIZE),
				to_sfixed(0.8723,1,L_SIZE),
				to_sfixed(0.8724,1,L_SIZE),
				to_sfixed(0.8725,1,L_SIZE),
				to_sfixed(0.8725,1,L_SIZE),
				to_sfixed(0.8726,1,L_SIZE),
				to_sfixed(0.8727,1,L_SIZE),
				to_sfixed(0.8728,1,L_SIZE),
				to_sfixed(0.8729,1,L_SIZE),
				to_sfixed(0.8730,1,L_SIZE),
				to_sfixed(0.8731,1,L_SIZE),
				to_sfixed(0.8732,1,L_SIZE),
				to_sfixed(0.8732,1,L_SIZE),
				to_sfixed(0.8733,1,L_SIZE),
				to_sfixed(0.8734,1,L_SIZE),
				to_sfixed(0.8735,1,L_SIZE),
				to_sfixed(0.8736,1,L_SIZE),
				to_sfixed(0.8737,1,L_SIZE),
				to_sfixed(0.8738,1,L_SIZE),
				to_sfixed(0.8738,1,L_SIZE),
				to_sfixed(0.8739,1,L_SIZE),
				to_sfixed(0.8740,1,L_SIZE),
				to_sfixed(0.8741,1,L_SIZE),
				to_sfixed(0.8742,1,L_SIZE),
				to_sfixed(0.8743,1,L_SIZE),
				to_sfixed(0.8744,1,L_SIZE),
				to_sfixed(0.8745,1,L_SIZE),
				to_sfixed(0.8745,1,L_SIZE),
				to_sfixed(0.8746,1,L_SIZE),
				to_sfixed(0.8747,1,L_SIZE),
				to_sfixed(0.8748,1,L_SIZE),
				to_sfixed(0.8749,1,L_SIZE),
				to_sfixed(0.8750,1,L_SIZE),
				to_sfixed(0.8751,1,L_SIZE),
				to_sfixed(0.8751,1,L_SIZE),
				to_sfixed(0.8752,1,L_SIZE),
				to_sfixed(0.8753,1,L_SIZE),
				to_sfixed(0.8754,1,L_SIZE),
				to_sfixed(0.8755,1,L_SIZE),
				to_sfixed(0.8756,1,L_SIZE),
				to_sfixed(0.8757,1,L_SIZE),
				to_sfixed(0.8757,1,L_SIZE),
				to_sfixed(0.8758,1,L_SIZE),
				to_sfixed(0.8759,1,L_SIZE),
				to_sfixed(0.8760,1,L_SIZE),
				to_sfixed(0.8761,1,L_SIZE),
				to_sfixed(0.8762,1,L_SIZE),
				to_sfixed(0.8762,1,L_SIZE),
				to_sfixed(0.8763,1,L_SIZE),
				to_sfixed(0.8764,1,L_SIZE),
				to_sfixed(0.8765,1,L_SIZE),
				to_sfixed(0.8766,1,L_SIZE),
				to_sfixed(0.8767,1,L_SIZE),
				to_sfixed(0.8768,1,L_SIZE),
				to_sfixed(0.8768,1,L_SIZE),
				to_sfixed(0.8769,1,L_SIZE),
				to_sfixed(0.8770,1,L_SIZE),
				to_sfixed(0.8771,1,L_SIZE),
				to_sfixed(0.8772,1,L_SIZE),
				to_sfixed(0.8773,1,L_SIZE),
				to_sfixed(0.8773,1,L_SIZE),
				to_sfixed(0.8774,1,L_SIZE),
				to_sfixed(0.8775,1,L_SIZE),
				to_sfixed(0.8776,1,L_SIZE),
				to_sfixed(0.8777,1,L_SIZE),
				to_sfixed(0.8778,1,L_SIZE),
				to_sfixed(0.8779,1,L_SIZE),
				to_sfixed(0.8779,1,L_SIZE),
				to_sfixed(0.8780,1,L_SIZE),
				to_sfixed(0.8781,1,L_SIZE),
				to_sfixed(0.8782,1,L_SIZE),
				to_sfixed(0.8783,1,L_SIZE),
				to_sfixed(0.8784,1,L_SIZE),
				to_sfixed(0.8784,1,L_SIZE),
				to_sfixed(0.8785,1,L_SIZE),
				to_sfixed(0.8786,1,L_SIZE),
				to_sfixed(0.8787,1,L_SIZE),
				to_sfixed(0.8788,1,L_SIZE),
				to_sfixed(0.8789,1,L_SIZE),
				to_sfixed(0.8789,1,L_SIZE),
				to_sfixed(0.8790,1,L_SIZE),
				to_sfixed(0.8791,1,L_SIZE),
				to_sfixed(0.8792,1,L_SIZE),
				to_sfixed(0.8793,1,L_SIZE),
				to_sfixed(0.8794,1,L_SIZE),
				to_sfixed(0.8794,1,L_SIZE),
				to_sfixed(0.8795,1,L_SIZE),
				to_sfixed(0.8796,1,L_SIZE),
				to_sfixed(0.8797,1,L_SIZE),
				to_sfixed(0.8798,1,L_SIZE),
				to_sfixed(0.8799,1,L_SIZE),
				to_sfixed(0.8799,1,L_SIZE),
				to_sfixed(0.8800,1,L_SIZE),
				to_sfixed(0.8801,1,L_SIZE),
				to_sfixed(0.8802,1,L_SIZE),
				to_sfixed(0.8803,1,L_SIZE),
				to_sfixed(0.8803,1,L_SIZE),
				to_sfixed(0.8804,1,L_SIZE),
				to_sfixed(0.8805,1,L_SIZE),
				to_sfixed(0.8806,1,L_SIZE),
				to_sfixed(0.8807,1,L_SIZE),
				to_sfixed(0.8808,1,L_SIZE),
				to_sfixed(0.8808,1,L_SIZE),
				to_sfixed(0.8809,1,L_SIZE),
				to_sfixed(0.8810,1,L_SIZE),
				to_sfixed(0.8811,1,L_SIZE),
				to_sfixed(0.8812,1,L_SIZE),
				to_sfixed(0.8813,1,L_SIZE),
				to_sfixed(0.8813,1,L_SIZE),
				to_sfixed(0.8814,1,L_SIZE),
				to_sfixed(0.8815,1,L_SIZE),
				to_sfixed(0.8816,1,L_SIZE),
				to_sfixed(0.8817,1,L_SIZE),
				to_sfixed(0.8817,1,L_SIZE),
				to_sfixed(0.8818,1,L_SIZE),
				to_sfixed(0.8819,1,L_SIZE),
				to_sfixed(0.8820,1,L_SIZE),
				to_sfixed(0.8821,1,L_SIZE),
				to_sfixed(0.8821,1,L_SIZE),
				to_sfixed(0.8822,1,L_SIZE),
				to_sfixed(0.8823,1,L_SIZE),
				to_sfixed(0.8824,1,L_SIZE),
				to_sfixed(0.8825,1,L_SIZE),
				to_sfixed(0.8826,1,L_SIZE),
				to_sfixed(0.8826,1,L_SIZE),
				to_sfixed(0.8827,1,L_SIZE),
				to_sfixed(0.8828,1,L_SIZE),
				to_sfixed(0.8829,1,L_SIZE),
				to_sfixed(0.8830,1,L_SIZE),
				to_sfixed(0.8830,1,L_SIZE),
				to_sfixed(0.8831,1,L_SIZE),
				to_sfixed(0.8832,1,L_SIZE),
				to_sfixed(0.8833,1,L_SIZE),
				to_sfixed(0.8834,1,L_SIZE),
				to_sfixed(0.8834,1,L_SIZE),
				to_sfixed(0.8835,1,L_SIZE),
				to_sfixed(0.8836,1,L_SIZE),
				to_sfixed(0.8837,1,L_SIZE),
				to_sfixed(0.8838,1,L_SIZE),
				to_sfixed(0.8838,1,L_SIZE),
				to_sfixed(0.8839,1,L_SIZE),
				to_sfixed(0.8840,1,L_SIZE),
				to_sfixed(0.8841,1,L_SIZE),
				to_sfixed(0.8842,1,L_SIZE),
				to_sfixed(0.8842,1,L_SIZE),
				to_sfixed(0.8843,1,L_SIZE),
				to_sfixed(0.8844,1,L_SIZE),
				to_sfixed(0.8845,1,L_SIZE),
				to_sfixed(0.8846,1,L_SIZE),
				to_sfixed(0.8846,1,L_SIZE),
				to_sfixed(0.8847,1,L_SIZE),
				to_sfixed(0.8848,1,L_SIZE),
				to_sfixed(0.8849,1,L_SIZE),
				to_sfixed(0.8850,1,L_SIZE),
				to_sfixed(0.8850,1,L_SIZE),
				to_sfixed(0.8851,1,L_SIZE),
				to_sfixed(0.8852,1,L_SIZE),
				to_sfixed(0.8853,1,L_SIZE),
				to_sfixed(0.8854,1,L_SIZE),
				to_sfixed(0.8854,1,L_SIZE),
				to_sfixed(0.8855,1,L_SIZE),
				to_sfixed(0.8856,1,L_SIZE),
				to_sfixed(0.8857,1,L_SIZE),
				to_sfixed(0.8858,1,L_SIZE),
				to_sfixed(0.8858,1,L_SIZE),
				to_sfixed(0.8859,1,L_SIZE),
				to_sfixed(0.8860,1,L_SIZE),
				to_sfixed(0.8861,1,L_SIZE),
				to_sfixed(0.8861,1,L_SIZE),
				to_sfixed(0.8862,1,L_SIZE),
				to_sfixed(0.8863,1,L_SIZE),
				to_sfixed(0.8864,1,L_SIZE),
				to_sfixed(0.8865,1,L_SIZE),
				to_sfixed(0.8865,1,L_SIZE),
				to_sfixed(0.8866,1,L_SIZE),
				to_sfixed(0.8867,1,L_SIZE),
				to_sfixed(0.8868,1,L_SIZE),
				to_sfixed(0.8869,1,L_SIZE),
				to_sfixed(0.8869,1,L_SIZE),
				to_sfixed(0.8870,1,L_SIZE),
				to_sfixed(0.8871,1,L_SIZE),
				to_sfixed(0.8872,1,L_SIZE),
				to_sfixed(0.8872,1,L_SIZE),
				to_sfixed(0.8873,1,L_SIZE),
				to_sfixed(0.8874,1,L_SIZE),
				to_sfixed(0.8875,1,L_SIZE),
				to_sfixed(0.8876,1,L_SIZE),
				to_sfixed(0.8876,1,L_SIZE),
				to_sfixed(0.8877,1,L_SIZE),
				to_sfixed(0.8878,1,L_SIZE),
				to_sfixed(0.8879,1,L_SIZE),
				to_sfixed(0.8879,1,L_SIZE),
				to_sfixed(0.8880,1,L_SIZE),
				to_sfixed(0.8881,1,L_SIZE),
				to_sfixed(0.8882,1,L_SIZE),
				to_sfixed(0.8883,1,L_SIZE),
				to_sfixed(0.8883,1,L_SIZE),
				to_sfixed(0.8884,1,L_SIZE),
				to_sfixed(0.8885,1,L_SIZE),
				to_sfixed(0.8886,1,L_SIZE),
				to_sfixed(0.8886,1,L_SIZE),
				to_sfixed(0.8887,1,L_SIZE),
				to_sfixed(0.8888,1,L_SIZE),
				to_sfixed(0.8889,1,L_SIZE),
				to_sfixed(0.8889,1,L_SIZE),
				to_sfixed(0.8890,1,L_SIZE),
				to_sfixed(0.8891,1,L_SIZE),
				to_sfixed(0.8892,1,L_SIZE),
				to_sfixed(0.8893,1,L_SIZE),
				to_sfixed(0.8893,1,L_SIZE),
				to_sfixed(0.8894,1,L_SIZE),
				to_sfixed(0.8895,1,L_SIZE),
				to_sfixed(0.8896,1,L_SIZE),
				to_sfixed(0.8896,1,L_SIZE),
				to_sfixed(0.8897,1,L_SIZE),
				to_sfixed(0.8898,1,L_SIZE),
				to_sfixed(0.8899,1,L_SIZE),
				to_sfixed(0.8899,1,L_SIZE),
				to_sfixed(0.8900,1,L_SIZE),
				to_sfixed(0.8901,1,L_SIZE),
				to_sfixed(0.8902,1,L_SIZE),
				to_sfixed(0.8902,1,L_SIZE),
				to_sfixed(0.8903,1,L_SIZE),
				to_sfixed(0.8904,1,L_SIZE),
				to_sfixed(0.8905,1,L_SIZE),
				to_sfixed(0.8905,1,L_SIZE),
				to_sfixed(0.8906,1,L_SIZE),
				to_sfixed(0.8907,1,L_SIZE),
				to_sfixed(0.8908,1,L_SIZE),
				to_sfixed(0.8908,1,L_SIZE),
				to_sfixed(0.8909,1,L_SIZE),
				to_sfixed(0.8910,1,L_SIZE),
				to_sfixed(0.8911,1,L_SIZE),
				to_sfixed(0.8912,1,L_SIZE),
				to_sfixed(0.8912,1,L_SIZE),
				to_sfixed(0.8913,1,L_SIZE),
				to_sfixed(0.8914,1,L_SIZE),
				to_sfixed(0.8915,1,L_SIZE),
				to_sfixed(0.8915,1,L_SIZE),
				to_sfixed(0.8916,1,L_SIZE),
				to_sfixed(0.8917,1,L_SIZE),
				to_sfixed(0.8918,1,L_SIZE),
				to_sfixed(0.8918,1,L_SIZE),
				to_sfixed(0.8919,1,L_SIZE),
				to_sfixed(0.8920,1,L_SIZE),
				to_sfixed(0.8921,1,L_SIZE),
				to_sfixed(0.8921,1,L_SIZE),
				to_sfixed(0.8922,1,L_SIZE),
				to_sfixed(0.8923,1,L_SIZE),
				to_sfixed(0.8924,1,L_SIZE),
				to_sfixed(0.8924,1,L_SIZE),
				to_sfixed(0.8925,1,L_SIZE),
				to_sfixed(0.8926,1,L_SIZE),
				to_sfixed(0.8926,1,L_SIZE),
				to_sfixed(0.8927,1,L_SIZE),
				to_sfixed(0.8928,1,L_SIZE),
				to_sfixed(0.8929,1,L_SIZE),
				to_sfixed(0.8929,1,L_SIZE),
				to_sfixed(0.8930,1,L_SIZE),
				to_sfixed(0.8931,1,L_SIZE),
				to_sfixed(0.8932,1,L_SIZE),
				to_sfixed(0.8932,1,L_SIZE),
				to_sfixed(0.8933,1,L_SIZE),
				to_sfixed(0.8934,1,L_SIZE),
				to_sfixed(0.8935,1,L_SIZE),
				to_sfixed(0.8935,1,L_SIZE),
				to_sfixed(0.8936,1,L_SIZE),
				to_sfixed(0.8937,1,L_SIZE),
				to_sfixed(0.8938,1,L_SIZE),
				to_sfixed(0.8938,1,L_SIZE),
				to_sfixed(0.8939,1,L_SIZE),
				to_sfixed(0.8940,1,L_SIZE),
				to_sfixed(0.8941,1,L_SIZE),
				to_sfixed(0.8941,1,L_SIZE),
				to_sfixed(0.8942,1,L_SIZE),
				to_sfixed(0.8943,1,L_SIZE),
				to_sfixed(0.8943,1,L_SIZE),
				to_sfixed(0.8944,1,L_SIZE),
				to_sfixed(0.8945,1,L_SIZE),
				to_sfixed(0.8946,1,L_SIZE),
				to_sfixed(0.8946,1,L_SIZE),
				to_sfixed(0.8947,1,L_SIZE),
				to_sfixed(0.8948,1,L_SIZE),
				to_sfixed(0.8949,1,L_SIZE),
				to_sfixed(0.8949,1,L_SIZE),
				to_sfixed(0.8950,1,L_SIZE),
				to_sfixed(0.8951,1,L_SIZE),
				to_sfixed(0.8952,1,L_SIZE),
				to_sfixed(0.8952,1,L_SIZE),
				to_sfixed(0.8953,1,L_SIZE),
				to_sfixed(0.8954,1,L_SIZE),
				to_sfixed(0.8954,1,L_SIZE),
				to_sfixed(0.8955,1,L_SIZE),
				to_sfixed(0.8956,1,L_SIZE),
				to_sfixed(0.8957,1,L_SIZE),
				to_sfixed(0.8957,1,L_SIZE),
				to_sfixed(0.8958,1,L_SIZE),
				to_sfixed(0.8959,1,L_SIZE),
				to_sfixed(0.8959,1,L_SIZE),
				to_sfixed(0.8960,1,L_SIZE),
				to_sfixed(0.8961,1,L_SIZE),
				to_sfixed(0.8962,1,L_SIZE),
				to_sfixed(0.8962,1,L_SIZE),
				to_sfixed(0.8963,1,L_SIZE),
				to_sfixed(0.8964,1,L_SIZE),
				to_sfixed(0.8965,1,L_SIZE),
				to_sfixed(0.8965,1,L_SIZE),
				to_sfixed(0.8966,1,L_SIZE),
				to_sfixed(0.8967,1,L_SIZE),
				to_sfixed(0.8967,1,L_SIZE),
				to_sfixed(0.8968,1,L_SIZE),
				to_sfixed(0.8969,1,L_SIZE),
				to_sfixed(0.8970,1,L_SIZE),
				to_sfixed(0.8970,1,L_SIZE),
				to_sfixed(0.8971,1,L_SIZE),
				to_sfixed(0.8972,1,L_SIZE),
				to_sfixed(0.8972,1,L_SIZE),
				to_sfixed(0.8973,1,L_SIZE),
				to_sfixed(0.8974,1,L_SIZE),
				to_sfixed(0.8975,1,L_SIZE),
				to_sfixed(0.8975,1,L_SIZE),
				to_sfixed(0.8976,1,L_SIZE),
				to_sfixed(0.8977,1,L_SIZE),
				to_sfixed(0.8977,1,L_SIZE),
				to_sfixed(0.8978,1,L_SIZE),
				to_sfixed(0.8979,1,L_SIZE),
				to_sfixed(0.8980,1,L_SIZE),
				to_sfixed(0.8980,1,L_SIZE),
				to_sfixed(0.8981,1,L_SIZE),
				to_sfixed(0.8982,1,L_SIZE),
				to_sfixed(0.8982,1,L_SIZE),
				to_sfixed(0.8983,1,L_SIZE),
				to_sfixed(0.8984,1,L_SIZE),
				to_sfixed(0.8984,1,L_SIZE),
				to_sfixed(0.8985,1,L_SIZE),
				to_sfixed(0.8986,1,L_SIZE),
				to_sfixed(0.8987,1,L_SIZE),
				to_sfixed(0.8987,1,L_SIZE),
				to_sfixed(0.8988,1,L_SIZE),
				to_sfixed(0.8989,1,L_SIZE),
				to_sfixed(0.8989,1,L_SIZE),
				to_sfixed(0.8990,1,L_SIZE),
				to_sfixed(0.8991,1,L_SIZE),
				to_sfixed(0.8992,1,L_SIZE),
				to_sfixed(0.8992,1,L_SIZE),
				to_sfixed(0.8993,1,L_SIZE),
				to_sfixed(0.8994,1,L_SIZE),
				to_sfixed(0.8994,1,L_SIZE),
				to_sfixed(0.8995,1,L_SIZE),
				to_sfixed(0.8996,1,L_SIZE),
				to_sfixed(0.8996,1,L_SIZE),
				to_sfixed(0.8997,1,L_SIZE),
				to_sfixed(0.8998,1,L_SIZE),
				to_sfixed(0.8999,1,L_SIZE),
				to_sfixed(0.8999,1,L_SIZE),
				to_sfixed(0.9000,1,L_SIZE),
				to_sfixed(0.9001,1,L_SIZE),
				to_sfixed(0.9001,1,L_SIZE),
				to_sfixed(0.9002,1,L_SIZE),
				to_sfixed(0.9003,1,L_SIZE),
				to_sfixed(0.9003,1,L_SIZE),
				to_sfixed(0.9004,1,L_SIZE),
				to_sfixed(0.9005,1,L_SIZE),
				to_sfixed(0.9005,1,L_SIZE),
				to_sfixed(0.9006,1,L_SIZE),
				to_sfixed(0.9007,1,L_SIZE),
				to_sfixed(0.9008,1,L_SIZE),
				to_sfixed(0.9008,1,L_SIZE),
				to_sfixed(0.9009,1,L_SIZE),
				to_sfixed(0.9010,1,L_SIZE),
				to_sfixed(0.9010,1,L_SIZE),
				to_sfixed(0.9011,1,L_SIZE),
				to_sfixed(0.9012,1,L_SIZE),
				to_sfixed(0.9012,1,L_SIZE),
				to_sfixed(0.9013,1,L_SIZE),
				to_sfixed(0.9014,1,L_SIZE),
				to_sfixed(0.9014,1,L_SIZE),
				to_sfixed(0.9015,1,L_SIZE),
				to_sfixed(0.9016,1,L_SIZE),
				to_sfixed(0.9016,1,L_SIZE),
				to_sfixed(0.9017,1,L_SIZE),
				to_sfixed(0.9018,1,L_SIZE),
				to_sfixed(0.9019,1,L_SIZE),
				to_sfixed(0.9019,1,L_SIZE),
				to_sfixed(0.9020,1,L_SIZE),
				to_sfixed(0.9021,1,L_SIZE),
				to_sfixed(0.9021,1,L_SIZE),
				to_sfixed(0.9022,1,L_SIZE),
				to_sfixed(0.9023,1,L_SIZE),
				to_sfixed(0.9023,1,L_SIZE),
				to_sfixed(0.9024,1,L_SIZE),
				to_sfixed(0.9025,1,L_SIZE),
				to_sfixed(0.9025,1,L_SIZE),
				to_sfixed(0.9026,1,L_SIZE),
				to_sfixed(0.9027,1,L_SIZE),
				to_sfixed(0.9027,1,L_SIZE),
				to_sfixed(0.9028,1,L_SIZE),
				to_sfixed(0.9029,1,L_SIZE),
				to_sfixed(0.9029,1,L_SIZE),
				to_sfixed(0.9030,1,L_SIZE),
				to_sfixed(0.9031,1,L_SIZE),
				to_sfixed(0.9031,1,L_SIZE),
				to_sfixed(0.9032,1,L_SIZE),
				to_sfixed(0.9033,1,L_SIZE),
				to_sfixed(0.9033,1,L_SIZE),
				to_sfixed(0.9034,1,L_SIZE),
				to_sfixed(0.9035,1,L_SIZE),
				to_sfixed(0.9035,1,L_SIZE),
				to_sfixed(0.9036,1,L_SIZE),
				to_sfixed(0.9037,1,L_SIZE),
				to_sfixed(0.9037,1,L_SIZE),
				to_sfixed(0.9038,1,L_SIZE),
				to_sfixed(0.9039,1,L_SIZE),
				to_sfixed(0.9039,1,L_SIZE),
				to_sfixed(0.9040,1,L_SIZE),
				to_sfixed(0.9041,1,L_SIZE),
				to_sfixed(0.9042,1,L_SIZE),
				to_sfixed(0.9042,1,L_SIZE),
				to_sfixed(0.9043,1,L_SIZE),
				to_sfixed(0.9044,1,L_SIZE),
				to_sfixed(0.9044,1,L_SIZE),
				to_sfixed(0.9045,1,L_SIZE),
				to_sfixed(0.9046,1,L_SIZE),
				to_sfixed(0.9046,1,L_SIZE),
				to_sfixed(0.9047,1,L_SIZE),
				to_sfixed(0.9048,1,L_SIZE),
				to_sfixed(0.9048,1,L_SIZE),
				to_sfixed(0.9049,1,L_SIZE),
				to_sfixed(0.9049,1,L_SIZE),
				to_sfixed(0.9050,1,L_SIZE),
				to_sfixed(0.9051,1,L_SIZE),
				to_sfixed(0.9051,1,L_SIZE),
				to_sfixed(0.9052,1,L_SIZE),
				to_sfixed(0.9053,1,L_SIZE),
				to_sfixed(0.9053,1,L_SIZE),
				to_sfixed(0.9054,1,L_SIZE),
				to_sfixed(0.9055,1,L_SIZE),
				to_sfixed(0.9055,1,L_SIZE),
				to_sfixed(0.9056,1,L_SIZE),
				to_sfixed(0.9057,1,L_SIZE),
				to_sfixed(0.9057,1,L_SIZE),
				to_sfixed(0.9058,1,L_SIZE),
				to_sfixed(0.9059,1,L_SIZE),
				to_sfixed(0.9059,1,L_SIZE),
				to_sfixed(0.9060,1,L_SIZE),
				to_sfixed(0.9061,1,L_SIZE),
				to_sfixed(0.9061,1,L_SIZE),
				to_sfixed(0.9062,1,L_SIZE),
				to_sfixed(0.9063,1,L_SIZE),
				to_sfixed(0.9063,1,L_SIZE),
				to_sfixed(0.9064,1,L_SIZE),
				to_sfixed(0.9065,1,L_SIZE),
				to_sfixed(0.9065,1,L_SIZE),
				to_sfixed(0.9066,1,L_SIZE),
				to_sfixed(0.9067,1,L_SIZE),
				to_sfixed(0.9067,1,L_SIZE),
				to_sfixed(0.9068,1,L_SIZE),
				to_sfixed(0.9069,1,L_SIZE),
				to_sfixed(0.9069,1,L_SIZE),
				to_sfixed(0.9070,1,L_SIZE),
				to_sfixed(0.9070,1,L_SIZE),
				to_sfixed(0.9071,1,L_SIZE),
				to_sfixed(0.9072,1,L_SIZE),
				to_sfixed(0.9072,1,L_SIZE),
				to_sfixed(0.9073,1,L_SIZE),
				to_sfixed(0.9074,1,L_SIZE),
				to_sfixed(0.9074,1,L_SIZE),
				to_sfixed(0.9075,1,L_SIZE),
				to_sfixed(0.9076,1,L_SIZE),
				to_sfixed(0.9076,1,L_SIZE),
				to_sfixed(0.9077,1,L_SIZE),
				to_sfixed(0.9078,1,L_SIZE),
				to_sfixed(0.9078,1,L_SIZE),
				to_sfixed(0.9079,1,L_SIZE),
				to_sfixed(0.9080,1,L_SIZE),
				to_sfixed(0.9080,1,L_SIZE),
				to_sfixed(0.9081,1,L_SIZE),
				to_sfixed(0.9081,1,L_SIZE),
				to_sfixed(0.9082,1,L_SIZE),
				to_sfixed(0.9083,1,L_SIZE),
				to_sfixed(0.9083,1,L_SIZE),
				to_sfixed(0.9084,1,L_SIZE),
				to_sfixed(0.9085,1,L_SIZE),
				to_sfixed(0.9085,1,L_SIZE),
				to_sfixed(0.9086,1,L_SIZE),
				to_sfixed(0.9087,1,L_SIZE),
				to_sfixed(0.9087,1,L_SIZE),
				to_sfixed(0.9088,1,L_SIZE),
				to_sfixed(0.9088,1,L_SIZE),
				to_sfixed(0.9089,1,L_SIZE),
				to_sfixed(0.9090,1,L_SIZE),
				to_sfixed(0.9090,1,L_SIZE),
				to_sfixed(0.9091,1,L_SIZE),
				to_sfixed(0.9092,1,L_SIZE),
				to_sfixed(0.9092,1,L_SIZE),
				to_sfixed(0.9093,1,L_SIZE),
				to_sfixed(0.9094,1,L_SIZE),
				to_sfixed(0.9094,1,L_SIZE),
				to_sfixed(0.9095,1,L_SIZE),
				to_sfixed(0.9095,1,L_SIZE),
				to_sfixed(0.9096,1,L_SIZE),
				to_sfixed(0.9097,1,L_SIZE),
				to_sfixed(0.9097,1,L_SIZE),
				to_sfixed(0.9098,1,L_SIZE),
				to_sfixed(0.9099,1,L_SIZE),
				to_sfixed(0.9099,1,L_SIZE),
				to_sfixed(0.9100,1,L_SIZE),
				to_sfixed(0.9101,1,L_SIZE),
				to_sfixed(0.9101,1,L_SIZE),
				to_sfixed(0.9102,1,L_SIZE),
				to_sfixed(0.9102,1,L_SIZE),
				to_sfixed(0.9103,1,L_SIZE),
				to_sfixed(0.9104,1,L_SIZE),
				to_sfixed(0.9104,1,L_SIZE),
				to_sfixed(0.9105,1,L_SIZE),
				to_sfixed(0.9106,1,L_SIZE),
				to_sfixed(0.9106,1,L_SIZE),
				to_sfixed(0.9107,1,L_SIZE),
				to_sfixed(0.9107,1,L_SIZE),
				to_sfixed(0.9108,1,L_SIZE),
				to_sfixed(0.9109,1,L_SIZE),
				to_sfixed(0.9109,1,L_SIZE),
				to_sfixed(0.9110,1,L_SIZE),
				to_sfixed(0.9111,1,L_SIZE),
				to_sfixed(0.9111,1,L_SIZE),
				to_sfixed(0.9112,1,L_SIZE),
				to_sfixed(0.9112,1,L_SIZE),
				to_sfixed(0.9113,1,L_SIZE),
				to_sfixed(0.9114,1,L_SIZE),
				to_sfixed(0.9114,1,L_SIZE),
				to_sfixed(0.9115,1,L_SIZE),
				to_sfixed(0.9116,1,L_SIZE),
				to_sfixed(0.9116,1,L_SIZE),
				to_sfixed(0.9117,1,L_SIZE),
				to_sfixed(0.9117,1,L_SIZE),
				to_sfixed(0.9118,1,L_SIZE),
				to_sfixed(0.9119,1,L_SIZE),
				to_sfixed(0.9119,1,L_SIZE),
				to_sfixed(0.9120,1,L_SIZE),
				to_sfixed(0.9120,1,L_SIZE),
				to_sfixed(0.9121,1,L_SIZE),
				to_sfixed(0.9122,1,L_SIZE),
				to_sfixed(0.9122,1,L_SIZE),
				to_sfixed(0.9123,1,L_SIZE),
				to_sfixed(0.9124,1,L_SIZE),
				to_sfixed(0.9124,1,L_SIZE),
				to_sfixed(0.9125,1,L_SIZE),
				to_sfixed(0.9125,1,L_SIZE),
				to_sfixed(0.9126,1,L_SIZE),
				to_sfixed(0.9127,1,L_SIZE),
				to_sfixed(0.9127,1,L_SIZE),
				to_sfixed(0.9128,1,L_SIZE),
				to_sfixed(0.9128,1,L_SIZE),
				to_sfixed(0.9129,1,L_SIZE),
				to_sfixed(0.9130,1,L_SIZE),
				to_sfixed(0.9130,1,L_SIZE),
				to_sfixed(0.9131,1,L_SIZE),
				to_sfixed(0.9131,1,L_SIZE),
				to_sfixed(0.9132,1,L_SIZE),
				to_sfixed(0.9133,1,L_SIZE),
				to_sfixed(0.9133,1,L_SIZE),
				to_sfixed(0.9134,1,L_SIZE),
				to_sfixed(0.9135,1,L_SIZE),
				to_sfixed(0.9135,1,L_SIZE),
				to_sfixed(0.9136,1,L_SIZE),
				to_sfixed(0.9136,1,L_SIZE),
				to_sfixed(0.9137,1,L_SIZE),
				to_sfixed(0.9138,1,L_SIZE),
				to_sfixed(0.9138,1,L_SIZE),
				to_sfixed(0.9139,1,L_SIZE),
				to_sfixed(0.9139,1,L_SIZE),
				to_sfixed(0.9140,1,L_SIZE),
				to_sfixed(0.9141,1,L_SIZE),
				to_sfixed(0.9141,1,L_SIZE),
				to_sfixed(0.9142,1,L_SIZE),
				to_sfixed(0.9142,1,L_SIZE),
				to_sfixed(0.9143,1,L_SIZE),
				to_sfixed(0.9144,1,L_SIZE),
				to_sfixed(0.9144,1,L_SIZE),
				to_sfixed(0.9145,1,L_SIZE),
				to_sfixed(0.9145,1,L_SIZE),
				to_sfixed(0.9146,1,L_SIZE),
				to_sfixed(0.9147,1,L_SIZE),
				to_sfixed(0.9147,1,L_SIZE),
				to_sfixed(0.9148,1,L_SIZE),
				to_sfixed(0.9148,1,L_SIZE),
				to_sfixed(0.9149,1,L_SIZE),
				to_sfixed(0.9150,1,L_SIZE),
				to_sfixed(0.9150,1,L_SIZE),
				to_sfixed(0.9151,1,L_SIZE),
				to_sfixed(0.9151,1,L_SIZE),
				to_sfixed(0.9152,1,L_SIZE),
				to_sfixed(0.9153,1,L_SIZE),
				to_sfixed(0.9153,1,L_SIZE),
				to_sfixed(0.9154,1,L_SIZE),
				to_sfixed(0.9154,1,L_SIZE),
				to_sfixed(0.9155,1,L_SIZE),
				to_sfixed(0.9155,1,L_SIZE),
				to_sfixed(0.9156,1,L_SIZE),
				to_sfixed(0.9157,1,L_SIZE),
				to_sfixed(0.9157,1,L_SIZE),
				to_sfixed(0.9158,1,L_SIZE),
				to_sfixed(0.9158,1,L_SIZE),
				to_sfixed(0.9159,1,L_SIZE),
				to_sfixed(0.9160,1,L_SIZE),
				to_sfixed(0.9160,1,L_SIZE),
				to_sfixed(0.9161,1,L_SIZE),
				to_sfixed(0.9161,1,L_SIZE),
				to_sfixed(0.9162,1,L_SIZE),
				to_sfixed(0.9163,1,L_SIZE),
				to_sfixed(0.9163,1,L_SIZE),
				to_sfixed(0.9164,1,L_SIZE),
				to_sfixed(0.9164,1,L_SIZE),
				to_sfixed(0.9165,1,L_SIZE),
				to_sfixed(0.9165,1,L_SIZE),
				to_sfixed(0.9166,1,L_SIZE),
				to_sfixed(0.9167,1,L_SIZE),
				to_sfixed(0.9167,1,L_SIZE),
				to_sfixed(0.9168,1,L_SIZE),
				to_sfixed(0.9168,1,L_SIZE),
				to_sfixed(0.9169,1,L_SIZE),
				to_sfixed(0.9170,1,L_SIZE),
				to_sfixed(0.9170,1,L_SIZE),
				to_sfixed(0.9171,1,L_SIZE),
				to_sfixed(0.9171,1,L_SIZE),
				to_sfixed(0.9172,1,L_SIZE),
				to_sfixed(0.9172,1,L_SIZE),
				to_sfixed(0.9173,1,L_SIZE),
				to_sfixed(0.9174,1,L_SIZE),
				to_sfixed(0.9174,1,L_SIZE),
				to_sfixed(0.9175,1,L_SIZE),
				to_sfixed(0.9175,1,L_SIZE),
				to_sfixed(0.9176,1,L_SIZE),
				to_sfixed(0.9177,1,L_SIZE),
				to_sfixed(0.9177,1,L_SIZE),
				to_sfixed(0.9178,1,L_SIZE),
				to_sfixed(0.9178,1,L_SIZE),
				to_sfixed(0.9179,1,L_SIZE),
				to_sfixed(0.9179,1,L_SIZE),
				to_sfixed(0.9180,1,L_SIZE),
				to_sfixed(0.9181,1,L_SIZE),
				to_sfixed(0.9181,1,L_SIZE),
				to_sfixed(0.9182,1,L_SIZE),
				to_sfixed(0.9182,1,L_SIZE),
				to_sfixed(0.9183,1,L_SIZE),
				to_sfixed(0.9183,1,L_SIZE),
				to_sfixed(0.9184,1,L_SIZE),
				to_sfixed(0.9185,1,L_SIZE),
				to_sfixed(0.9185,1,L_SIZE),
				to_sfixed(0.9186,1,L_SIZE),
				to_sfixed(0.9186,1,L_SIZE),
				to_sfixed(0.9187,1,L_SIZE),
				to_sfixed(0.9187,1,L_SIZE),
				to_sfixed(0.9188,1,L_SIZE),
				to_sfixed(0.9189,1,L_SIZE),
				to_sfixed(0.9189,1,L_SIZE),
				to_sfixed(0.9190,1,L_SIZE),
				to_sfixed(0.9190,1,L_SIZE),
				to_sfixed(0.9191,1,L_SIZE),
				to_sfixed(0.9191,1,L_SIZE),
				to_sfixed(0.9192,1,L_SIZE),
				to_sfixed(0.9193,1,L_SIZE),
				to_sfixed(0.9193,1,L_SIZE),
				to_sfixed(0.9194,1,L_SIZE),
				to_sfixed(0.9194,1,L_SIZE),
				to_sfixed(0.9195,1,L_SIZE),
				to_sfixed(0.9195,1,L_SIZE),
				to_sfixed(0.9196,1,L_SIZE),
				to_sfixed(0.9197,1,L_SIZE),
				to_sfixed(0.9197,1,L_SIZE),
				to_sfixed(0.9198,1,L_SIZE),
				to_sfixed(0.9198,1,L_SIZE),
				to_sfixed(0.9199,1,L_SIZE),
				to_sfixed(0.9199,1,L_SIZE),
				to_sfixed(0.9200,1,L_SIZE),
				to_sfixed(0.9201,1,L_SIZE),
				to_sfixed(0.9201,1,L_SIZE),
				to_sfixed(0.9202,1,L_SIZE),
				to_sfixed(0.9202,1,L_SIZE),
				to_sfixed(0.9203,1,L_SIZE),
				to_sfixed(0.9203,1,L_SIZE),
				to_sfixed(0.9204,1,L_SIZE),
				to_sfixed(0.9204,1,L_SIZE),
				to_sfixed(0.9205,1,L_SIZE),
				to_sfixed(0.9206,1,L_SIZE),
				to_sfixed(0.9206,1,L_SIZE),
				to_sfixed(0.9207,1,L_SIZE),
				to_sfixed(0.9207,1,L_SIZE),
				to_sfixed(0.9208,1,L_SIZE),
				to_sfixed(0.9208,1,L_SIZE),
				to_sfixed(0.9209,1,L_SIZE),
				to_sfixed(0.9209,1,L_SIZE),
				to_sfixed(0.9210,1,L_SIZE),
				to_sfixed(0.9211,1,L_SIZE),
				to_sfixed(0.9211,1,L_SIZE),
				to_sfixed(0.9212,1,L_SIZE),
				to_sfixed(0.9212,1,L_SIZE),
				to_sfixed(0.9213,1,L_SIZE),
				to_sfixed(0.9213,1,L_SIZE),
				to_sfixed(0.9214,1,L_SIZE),
				to_sfixed(0.9214,1,L_SIZE),
				to_sfixed(0.9215,1,L_SIZE),
				to_sfixed(0.9216,1,L_SIZE),
				to_sfixed(0.9216,1,L_SIZE),
				to_sfixed(0.9217,1,L_SIZE),
				to_sfixed(0.9217,1,L_SIZE),
				to_sfixed(0.9218,1,L_SIZE),
				to_sfixed(0.9218,1,L_SIZE),
				to_sfixed(0.9219,1,L_SIZE),
				to_sfixed(0.9219,1,L_SIZE),
				to_sfixed(0.9220,1,L_SIZE),
				to_sfixed(0.9220,1,L_SIZE),
				to_sfixed(0.9221,1,L_SIZE),
				to_sfixed(0.9222,1,L_SIZE),
				to_sfixed(0.9222,1,L_SIZE),
				to_sfixed(0.9223,1,L_SIZE),
				to_sfixed(0.9223,1,L_SIZE),
				to_sfixed(0.9224,1,L_SIZE),
				to_sfixed(0.9224,1,L_SIZE),
				to_sfixed(0.9225,1,L_SIZE),
				to_sfixed(0.9225,1,L_SIZE),
				to_sfixed(0.9226,1,L_SIZE),
				to_sfixed(0.9227,1,L_SIZE),
				to_sfixed(0.9227,1,L_SIZE),
				to_sfixed(0.9228,1,L_SIZE),
				to_sfixed(0.9228,1,L_SIZE),
				to_sfixed(0.9229,1,L_SIZE),
				to_sfixed(0.9229,1,L_SIZE),
				to_sfixed(0.9230,1,L_SIZE),
				to_sfixed(0.9230,1,L_SIZE),
				to_sfixed(0.9231,1,L_SIZE),
				to_sfixed(0.9231,1,L_SIZE),
				to_sfixed(0.9232,1,L_SIZE),
				to_sfixed(0.9232,1,L_SIZE),
				to_sfixed(0.9233,1,L_SIZE),
				to_sfixed(0.9234,1,L_SIZE),
				to_sfixed(0.9234,1,L_SIZE),
				to_sfixed(0.9235,1,L_SIZE),
				to_sfixed(0.9235,1,L_SIZE),
				to_sfixed(0.9236,1,L_SIZE),
				to_sfixed(0.9236,1,L_SIZE),
				to_sfixed(0.9237,1,L_SIZE),
				to_sfixed(0.9237,1,L_SIZE),
				to_sfixed(0.9238,1,L_SIZE),
				to_sfixed(0.9238,1,L_SIZE),
				to_sfixed(0.9239,1,L_SIZE),
				to_sfixed(0.9239,1,L_SIZE),
				to_sfixed(0.9240,1,L_SIZE),
				to_sfixed(0.9241,1,L_SIZE),
				to_sfixed(0.9241,1,L_SIZE),
				to_sfixed(0.9242,1,L_SIZE),
				to_sfixed(0.9242,1,L_SIZE),
				to_sfixed(0.9243,1,L_SIZE),
				to_sfixed(0.9243,1,L_SIZE),
				to_sfixed(0.9244,1,L_SIZE),
				to_sfixed(0.9244,1,L_SIZE),
				to_sfixed(0.9245,1,L_SIZE),
				to_sfixed(0.9245,1,L_SIZE),
				to_sfixed(0.9246,1,L_SIZE),
				to_sfixed(0.9246,1,L_SIZE),
				to_sfixed(0.9247,1,L_SIZE),
				to_sfixed(0.9247,1,L_SIZE),
				to_sfixed(0.9248,1,L_SIZE),
				to_sfixed(0.9249,1,L_SIZE),
				to_sfixed(0.9249,1,L_SIZE),
				to_sfixed(0.9250,1,L_SIZE),
				to_sfixed(0.9250,1,L_SIZE),
				to_sfixed(0.9251,1,L_SIZE),
				to_sfixed(0.9251,1,L_SIZE),
				to_sfixed(0.9252,1,L_SIZE),
				to_sfixed(0.9252,1,L_SIZE),
				to_sfixed(0.9253,1,L_SIZE),
				to_sfixed(0.9253,1,L_SIZE),
				to_sfixed(0.9254,1,L_SIZE),
				to_sfixed(0.9254,1,L_SIZE),
				to_sfixed(0.9255,1,L_SIZE),
				to_sfixed(0.9255,1,L_SIZE),
				to_sfixed(0.9256,1,L_SIZE),
				to_sfixed(0.9256,1,L_SIZE),
				to_sfixed(0.9257,1,L_SIZE),
				to_sfixed(0.9257,1,L_SIZE),
				to_sfixed(0.9258,1,L_SIZE),
				to_sfixed(0.9259,1,L_SIZE),
				to_sfixed(0.9259,1,L_SIZE),
				to_sfixed(0.9260,1,L_SIZE),
				to_sfixed(0.9260,1,L_SIZE),
				to_sfixed(0.9261,1,L_SIZE),
				to_sfixed(0.9261,1,L_SIZE),
				to_sfixed(0.9262,1,L_SIZE),
				to_sfixed(0.9262,1,L_SIZE),
				to_sfixed(0.9263,1,L_SIZE),
				to_sfixed(0.9263,1,L_SIZE),
				to_sfixed(0.9264,1,L_SIZE),
				to_sfixed(0.9264,1,L_SIZE),
				to_sfixed(0.9265,1,L_SIZE),
				to_sfixed(0.9265,1,L_SIZE),
				to_sfixed(0.9266,1,L_SIZE),
				to_sfixed(0.9266,1,L_SIZE),
				to_sfixed(0.9267,1,L_SIZE),
				to_sfixed(0.9267,1,L_SIZE),
				to_sfixed(0.9268,1,L_SIZE),
				to_sfixed(0.9268,1,L_SIZE),
				to_sfixed(0.9269,1,L_SIZE),
				to_sfixed(0.9269,1,L_SIZE),
				to_sfixed(0.9270,1,L_SIZE),
				to_sfixed(0.9270,1,L_SIZE),
				to_sfixed(0.9271,1,L_SIZE),
				to_sfixed(0.9271,1,L_SIZE),
				to_sfixed(0.9272,1,L_SIZE),
				to_sfixed(0.9273,1,L_SIZE),
				to_sfixed(0.9273,1,L_SIZE),
				to_sfixed(0.9274,1,L_SIZE),
				to_sfixed(0.9274,1,L_SIZE),
				to_sfixed(0.9275,1,L_SIZE),
				to_sfixed(0.9275,1,L_SIZE),
				to_sfixed(0.9276,1,L_SIZE),
				to_sfixed(0.9276,1,L_SIZE),
				to_sfixed(0.9277,1,L_SIZE),
				to_sfixed(0.9277,1,L_SIZE),
				to_sfixed(0.9278,1,L_SIZE),
				to_sfixed(0.9278,1,L_SIZE),
				to_sfixed(0.9279,1,L_SIZE),
				to_sfixed(0.9279,1,L_SIZE),
				to_sfixed(0.9280,1,L_SIZE),
				to_sfixed(0.9280,1,L_SIZE),
				to_sfixed(0.9281,1,L_SIZE),
				to_sfixed(0.9281,1,L_SIZE),
				to_sfixed(0.9282,1,L_SIZE),
				to_sfixed(0.9282,1,L_SIZE),
				to_sfixed(0.9283,1,L_SIZE),
				to_sfixed(0.9283,1,L_SIZE),
				to_sfixed(0.9284,1,L_SIZE),
				to_sfixed(0.9284,1,L_SIZE),
				to_sfixed(0.9285,1,L_SIZE),
				to_sfixed(0.9285,1,L_SIZE),
				to_sfixed(0.9286,1,L_SIZE),
				to_sfixed(0.9286,1,L_SIZE),
				to_sfixed(0.9287,1,L_SIZE),
				to_sfixed(0.9287,1,L_SIZE),
				to_sfixed(0.9288,1,L_SIZE),
				to_sfixed(0.9288,1,L_SIZE),
				to_sfixed(0.9289,1,L_SIZE),
				to_sfixed(0.9289,1,L_SIZE),
				to_sfixed(0.9290,1,L_SIZE),
				to_sfixed(0.9290,1,L_SIZE),
				to_sfixed(0.9291,1,L_SIZE),
				to_sfixed(0.9291,1,L_SIZE),
				to_sfixed(0.9292,1,L_SIZE),
				to_sfixed(0.9292,1,L_SIZE),
				to_sfixed(0.9293,1,L_SIZE),
				to_sfixed(0.9293,1,L_SIZE),
				to_sfixed(0.9294,1,L_SIZE),
				to_sfixed(0.9294,1,L_SIZE),
				to_sfixed(0.9295,1,L_SIZE),
				to_sfixed(0.9295,1,L_SIZE),
				to_sfixed(0.9296,1,L_SIZE),
				to_sfixed(0.9296,1,L_SIZE),
				to_sfixed(0.9297,1,L_SIZE),
				to_sfixed(0.9297,1,L_SIZE),
				to_sfixed(0.9298,1,L_SIZE),
				to_sfixed(0.9298,1,L_SIZE),
				to_sfixed(0.9299,1,L_SIZE),
				to_sfixed(0.9299,1,L_SIZE),
				to_sfixed(0.9300,1,L_SIZE),
				to_sfixed(0.9300,1,L_SIZE),
				to_sfixed(0.9301,1,L_SIZE),
				to_sfixed(0.9301,1,L_SIZE),
				to_sfixed(0.9302,1,L_SIZE),
				to_sfixed(0.9302,1,L_SIZE),
				to_sfixed(0.9303,1,L_SIZE),
				to_sfixed(0.9303,1,L_SIZE),
				to_sfixed(0.9304,1,L_SIZE),
				to_sfixed(0.9304,1,L_SIZE),
				to_sfixed(0.9305,1,L_SIZE),
				to_sfixed(0.9305,1,L_SIZE),
				to_sfixed(0.9306,1,L_SIZE),
				to_sfixed(0.9306,1,L_SIZE),
				to_sfixed(0.9307,1,L_SIZE),
				to_sfixed(0.9307,1,L_SIZE),
				to_sfixed(0.9308,1,L_SIZE),
				to_sfixed(0.9308,1,L_SIZE),
				to_sfixed(0.9309,1,L_SIZE),
				to_sfixed(0.9309,1,L_SIZE),
				to_sfixed(0.9310,1,L_SIZE),
				to_sfixed(0.9310,1,L_SIZE),
				to_sfixed(0.9311,1,L_SIZE),
				to_sfixed(0.9311,1,L_SIZE),
				to_sfixed(0.9312,1,L_SIZE),
				to_sfixed(0.9312,1,L_SIZE),
				to_sfixed(0.9313,1,L_SIZE),
				to_sfixed(0.9313,1,L_SIZE),
				to_sfixed(0.9313,1,L_SIZE),
				to_sfixed(0.9314,1,L_SIZE),
				to_sfixed(0.9314,1,L_SIZE),
				to_sfixed(0.9315,1,L_SIZE),
				to_sfixed(0.9315,1,L_SIZE),
				to_sfixed(0.9316,1,L_SIZE),
				to_sfixed(0.9316,1,L_SIZE),
				to_sfixed(0.9317,1,L_SIZE),
				to_sfixed(0.9317,1,L_SIZE),
				to_sfixed(0.9318,1,L_SIZE),
				to_sfixed(0.9318,1,L_SIZE),
				to_sfixed(0.9319,1,L_SIZE),
				to_sfixed(0.9319,1,L_SIZE),
				to_sfixed(0.9320,1,L_SIZE),
				to_sfixed(0.9320,1,L_SIZE),
				to_sfixed(0.9321,1,L_SIZE),
				to_sfixed(0.9321,1,L_SIZE),
				to_sfixed(0.9322,1,L_SIZE),
				to_sfixed(0.9322,1,L_SIZE),
				to_sfixed(0.9323,1,L_SIZE),
				to_sfixed(0.9323,1,L_SIZE),
				to_sfixed(0.9324,1,L_SIZE),
				to_sfixed(0.9324,1,L_SIZE),
				to_sfixed(0.9325,1,L_SIZE),
				to_sfixed(0.9325,1,L_SIZE),
				to_sfixed(0.9326,1,L_SIZE),
				to_sfixed(0.9326,1,L_SIZE),
				to_sfixed(0.9326,1,L_SIZE),
				to_sfixed(0.9327,1,L_SIZE),
				to_sfixed(0.9327,1,L_SIZE),
				to_sfixed(0.9328,1,L_SIZE),
				to_sfixed(0.9328,1,L_SIZE),
				to_sfixed(0.9329,1,L_SIZE),
				to_sfixed(0.9329,1,L_SIZE),
				to_sfixed(0.9330,1,L_SIZE),
				to_sfixed(0.9330,1,L_SIZE),
				to_sfixed(0.9331,1,L_SIZE),
				to_sfixed(0.9331,1,L_SIZE),
				to_sfixed(0.9332,1,L_SIZE),
				to_sfixed(0.9332,1,L_SIZE),
				to_sfixed(0.9333,1,L_SIZE),
				to_sfixed(0.9333,1,L_SIZE),
				to_sfixed(0.9334,1,L_SIZE),
				to_sfixed(0.9334,1,L_SIZE),
				to_sfixed(0.9335,1,L_SIZE),
				to_sfixed(0.9335,1,L_SIZE),
				to_sfixed(0.9335,1,L_SIZE),
				to_sfixed(0.9336,1,L_SIZE),
				to_sfixed(0.9336,1,L_SIZE),
				to_sfixed(0.9337,1,L_SIZE),
				to_sfixed(0.9337,1,L_SIZE),
				to_sfixed(0.9338,1,L_SIZE),
				to_sfixed(0.9338,1,L_SIZE),
				to_sfixed(0.9339,1,L_SIZE),
				to_sfixed(0.9339,1,L_SIZE),
				to_sfixed(0.9340,1,L_SIZE),
				to_sfixed(0.9340,1,L_SIZE),
				to_sfixed(0.9341,1,L_SIZE),
				to_sfixed(0.9341,1,L_SIZE),
				to_sfixed(0.9342,1,L_SIZE),
				to_sfixed(0.9342,1,L_SIZE),
				to_sfixed(0.9342,1,L_SIZE),
				to_sfixed(0.9343,1,L_SIZE),
				to_sfixed(0.9343,1,L_SIZE),
				to_sfixed(0.9344,1,L_SIZE),
				to_sfixed(0.9344,1,L_SIZE),
				to_sfixed(0.9345,1,L_SIZE),
				to_sfixed(0.9345,1,L_SIZE),
				to_sfixed(0.9346,1,L_SIZE),
				to_sfixed(0.9346,1,L_SIZE),
				to_sfixed(0.9347,1,L_SIZE),
				to_sfixed(0.9347,1,L_SIZE),
				to_sfixed(0.9348,1,L_SIZE),
				to_sfixed(0.9348,1,L_SIZE),
				to_sfixed(0.9349,1,L_SIZE),
				to_sfixed(0.9349,1,L_SIZE),
				to_sfixed(0.9349,1,L_SIZE),
				to_sfixed(0.9350,1,L_SIZE),
				to_sfixed(0.9350,1,L_SIZE),
				to_sfixed(0.9351,1,L_SIZE),
				to_sfixed(0.9351,1,L_SIZE),
				to_sfixed(0.9352,1,L_SIZE),
				to_sfixed(0.9352,1,L_SIZE),
				to_sfixed(0.9353,1,L_SIZE),
				to_sfixed(0.9353,1,L_SIZE),
				to_sfixed(0.9354,1,L_SIZE),
				to_sfixed(0.9354,1,L_SIZE),
				to_sfixed(0.9354,1,L_SIZE),
				to_sfixed(0.9355,1,L_SIZE),
				to_sfixed(0.9355,1,L_SIZE),
				to_sfixed(0.9356,1,L_SIZE),
				to_sfixed(0.9356,1,L_SIZE),
				to_sfixed(0.9357,1,L_SIZE),
				to_sfixed(0.9357,1,L_SIZE),
				to_sfixed(0.9358,1,L_SIZE),
				to_sfixed(0.9358,1,L_SIZE),
				to_sfixed(0.9359,1,L_SIZE),
				to_sfixed(0.9359,1,L_SIZE),
				to_sfixed(0.9360,1,L_SIZE),
				to_sfixed(0.9360,1,L_SIZE),
				to_sfixed(0.9360,1,L_SIZE),
				to_sfixed(0.9361,1,L_SIZE),
				to_sfixed(0.9361,1,L_SIZE),
				to_sfixed(0.9362,1,L_SIZE),
				to_sfixed(0.9362,1,L_SIZE),
				to_sfixed(0.9363,1,L_SIZE),
				to_sfixed(0.9363,1,L_SIZE),
				to_sfixed(0.9364,1,L_SIZE),
				to_sfixed(0.9364,1,L_SIZE),
				to_sfixed(0.9364,1,L_SIZE),
				to_sfixed(0.9365,1,L_SIZE),
				to_sfixed(0.9365,1,L_SIZE),
				to_sfixed(0.9366,1,L_SIZE),
				to_sfixed(0.9366,1,L_SIZE),
				to_sfixed(0.9367,1,L_SIZE),
				to_sfixed(0.9367,1,L_SIZE),
				to_sfixed(0.9368,1,L_SIZE),
				to_sfixed(0.9368,1,L_SIZE),
				to_sfixed(0.9369,1,L_SIZE),
				to_sfixed(0.9369,1,L_SIZE),
				to_sfixed(0.9369,1,L_SIZE),
				to_sfixed(0.9370,1,L_SIZE),
				to_sfixed(0.9370,1,L_SIZE),
				to_sfixed(0.9371,1,L_SIZE),
				to_sfixed(0.9371,1,L_SIZE),
				to_sfixed(0.9372,1,L_SIZE),
				to_sfixed(0.9372,1,L_SIZE),
				to_sfixed(0.9373,1,L_SIZE),
				to_sfixed(0.9373,1,L_SIZE),
				to_sfixed(0.9373,1,L_SIZE),
				to_sfixed(0.9374,1,L_SIZE),
				to_sfixed(0.9374,1,L_SIZE),
				to_sfixed(0.9375,1,L_SIZE),
				to_sfixed(0.9375,1,L_SIZE),
				to_sfixed(0.9376,1,L_SIZE),
				to_sfixed(0.9376,1,L_SIZE),
				to_sfixed(0.9377,1,L_SIZE),
				to_sfixed(0.9377,1,L_SIZE),
				to_sfixed(0.9377,1,L_SIZE),
				to_sfixed(0.9378,1,L_SIZE),
				to_sfixed(0.9378,1,L_SIZE),
				to_sfixed(0.9379,1,L_SIZE),
				to_sfixed(0.9379,1,L_SIZE),
				to_sfixed(0.9380,1,L_SIZE),
				to_sfixed(0.9380,1,L_SIZE),
				to_sfixed(0.9381,1,L_SIZE),
				to_sfixed(0.9381,1,L_SIZE),
				to_sfixed(0.9381,1,L_SIZE),
				to_sfixed(0.9382,1,L_SIZE),
				to_sfixed(0.9382,1,L_SIZE),
				to_sfixed(0.9383,1,L_SIZE),
				to_sfixed(0.9383,1,L_SIZE),
				to_sfixed(0.9384,1,L_SIZE),
				to_sfixed(0.9384,1,L_SIZE),
				to_sfixed(0.9384,1,L_SIZE),
				to_sfixed(0.9385,1,L_SIZE),
				to_sfixed(0.9385,1,L_SIZE),
				to_sfixed(0.9386,1,L_SIZE),
				to_sfixed(0.9386,1,L_SIZE),
				to_sfixed(0.9387,1,L_SIZE),
				to_sfixed(0.9387,1,L_SIZE),
				to_sfixed(0.9387,1,L_SIZE),
				to_sfixed(0.9388,1,L_SIZE),
				to_sfixed(0.9388,1,L_SIZE),
				to_sfixed(0.9389,1,L_SIZE),
				to_sfixed(0.9389,1,L_SIZE),
				to_sfixed(0.9390,1,L_SIZE),
				to_sfixed(0.9390,1,L_SIZE),
				to_sfixed(0.9391,1,L_SIZE),
				to_sfixed(0.9391,1,L_SIZE),
				to_sfixed(0.9391,1,L_SIZE),
				to_sfixed(0.9392,1,L_SIZE),
				to_sfixed(0.9392,1,L_SIZE),
				to_sfixed(0.9393,1,L_SIZE),
				to_sfixed(0.9393,1,L_SIZE),
				to_sfixed(0.9394,1,L_SIZE),
				to_sfixed(0.9394,1,L_SIZE),
				to_sfixed(0.9394,1,L_SIZE),
				to_sfixed(0.9395,1,L_SIZE),
				to_sfixed(0.9395,1,L_SIZE),
				to_sfixed(0.9396,1,L_SIZE),
				to_sfixed(0.9396,1,L_SIZE),
				to_sfixed(0.9397,1,L_SIZE),
				to_sfixed(0.9397,1,L_SIZE),
				to_sfixed(0.9397,1,L_SIZE),
				to_sfixed(0.9398,1,L_SIZE),
				to_sfixed(0.9398,1,L_SIZE),
				to_sfixed(0.9399,1,L_SIZE),
				to_sfixed(0.9399,1,L_SIZE),
				to_sfixed(0.9400,1,L_SIZE),
				to_sfixed(0.9400,1,L_SIZE),
				to_sfixed(0.9400,1,L_SIZE),
				to_sfixed(0.9401,1,L_SIZE),
				to_sfixed(0.9401,1,L_SIZE),
				to_sfixed(0.9402,1,L_SIZE),
				to_sfixed(0.9402,1,L_SIZE),
				to_sfixed(0.9403,1,L_SIZE),
				to_sfixed(0.9403,1,L_SIZE),
				to_sfixed(0.9403,1,L_SIZE),
				to_sfixed(0.9404,1,L_SIZE),
				to_sfixed(0.9404,1,L_SIZE),
				to_sfixed(0.9405,1,L_SIZE),
				to_sfixed(0.9405,1,L_SIZE),
				to_sfixed(0.9406,1,L_SIZE),
				to_sfixed(0.9406,1,L_SIZE),
				to_sfixed(0.9406,1,L_SIZE),
				to_sfixed(0.9407,1,L_SIZE),
				to_sfixed(0.9407,1,L_SIZE),
				to_sfixed(0.9408,1,L_SIZE),
				to_sfixed(0.9408,1,L_SIZE),
				to_sfixed(0.9408,1,L_SIZE),
				to_sfixed(0.9409,1,L_SIZE),
				to_sfixed(0.9409,1,L_SIZE),
				to_sfixed(0.9410,1,L_SIZE),
				to_sfixed(0.9410,1,L_SIZE),
				to_sfixed(0.9411,1,L_SIZE),
				to_sfixed(0.9411,1,L_SIZE),
				to_sfixed(0.9411,1,L_SIZE),
				to_sfixed(0.9412,1,L_SIZE),
				to_sfixed(0.9412,1,L_SIZE),
				to_sfixed(0.9413,1,L_SIZE),
				to_sfixed(0.9413,1,L_SIZE),
				to_sfixed(0.9413,1,L_SIZE),
				to_sfixed(0.9414,1,L_SIZE),
				to_sfixed(0.9414,1,L_SIZE),
				to_sfixed(0.9415,1,L_SIZE),
				to_sfixed(0.9415,1,L_SIZE),
				to_sfixed(0.9416,1,L_SIZE),
				to_sfixed(0.9416,1,L_SIZE),
				to_sfixed(0.9416,1,L_SIZE),
				to_sfixed(0.9417,1,L_SIZE),
				to_sfixed(0.9417,1,L_SIZE),
				to_sfixed(0.9418,1,L_SIZE),
				to_sfixed(0.9418,1,L_SIZE),
				to_sfixed(0.9418,1,L_SIZE),
				to_sfixed(0.9419,1,L_SIZE),
				to_sfixed(0.9419,1,L_SIZE),
				to_sfixed(0.9420,1,L_SIZE),
				to_sfixed(0.9420,1,L_SIZE),
				to_sfixed(0.9421,1,L_SIZE),
				to_sfixed(0.9421,1,L_SIZE),
				to_sfixed(0.9421,1,L_SIZE),
				to_sfixed(0.9422,1,L_SIZE),
				to_sfixed(0.9422,1,L_SIZE),
				to_sfixed(0.9423,1,L_SIZE),
				to_sfixed(0.9423,1,L_SIZE),
				to_sfixed(0.9423,1,L_SIZE),
				to_sfixed(0.9424,1,L_SIZE),
				to_sfixed(0.9424,1,L_SIZE),
				to_sfixed(0.9425,1,L_SIZE),
				to_sfixed(0.9425,1,L_SIZE),
				to_sfixed(0.9425,1,L_SIZE),
				to_sfixed(0.9426,1,L_SIZE),
				to_sfixed(0.9426,1,L_SIZE),
				to_sfixed(0.9427,1,L_SIZE),
				to_sfixed(0.9427,1,L_SIZE),
				to_sfixed(0.9427,1,L_SIZE),
				to_sfixed(0.9428,1,L_SIZE),
				to_sfixed(0.9428,1,L_SIZE),
				to_sfixed(0.9429,1,L_SIZE),
				to_sfixed(0.9429,1,L_SIZE),
				to_sfixed(0.9430,1,L_SIZE),
				to_sfixed(0.9430,1,L_SIZE),
				to_sfixed(0.9430,1,L_SIZE),
				to_sfixed(0.9431,1,L_SIZE),
				to_sfixed(0.9431,1,L_SIZE),
				to_sfixed(0.9432,1,L_SIZE),
				to_sfixed(0.9432,1,L_SIZE),
				to_sfixed(0.9432,1,L_SIZE),
				to_sfixed(0.9433,1,L_SIZE),
				to_sfixed(0.9433,1,L_SIZE),
				to_sfixed(0.9434,1,L_SIZE),
				to_sfixed(0.9434,1,L_SIZE),
				to_sfixed(0.9434,1,L_SIZE),
				to_sfixed(0.9435,1,L_SIZE),
				to_sfixed(0.9435,1,L_SIZE),
				to_sfixed(0.9436,1,L_SIZE),
				to_sfixed(0.9436,1,L_SIZE),
				to_sfixed(0.9436,1,L_SIZE),
				to_sfixed(0.9437,1,L_SIZE),
				to_sfixed(0.9437,1,L_SIZE),
				to_sfixed(0.9438,1,L_SIZE),
				to_sfixed(0.9438,1,L_SIZE),
				to_sfixed(0.9438,1,L_SIZE),
				to_sfixed(0.9439,1,L_SIZE),
				to_sfixed(0.9439,1,L_SIZE),
				to_sfixed(0.9440,1,L_SIZE),
				to_sfixed(0.9440,1,L_SIZE),
				to_sfixed(0.9440,1,L_SIZE),
				to_sfixed(0.9441,1,L_SIZE),
				to_sfixed(0.9441,1,L_SIZE),
				to_sfixed(0.9442,1,L_SIZE),
				to_sfixed(0.9442,1,L_SIZE),
				to_sfixed(0.9442,1,L_SIZE),
				to_sfixed(0.9443,1,L_SIZE),
				to_sfixed(0.9443,1,L_SIZE),
				to_sfixed(0.9444,1,L_SIZE),
				to_sfixed(0.9444,1,L_SIZE),
				to_sfixed(0.9444,1,L_SIZE),
				to_sfixed(0.9445,1,L_SIZE),
				to_sfixed(0.9445,1,L_SIZE),
				to_sfixed(0.9446,1,L_SIZE),
				to_sfixed(0.9446,1,L_SIZE),
				to_sfixed(0.9446,1,L_SIZE),
				to_sfixed(0.9447,1,L_SIZE),
				to_sfixed(0.9447,1,L_SIZE),
				to_sfixed(0.9448,1,L_SIZE),
				to_sfixed(0.9448,1,L_SIZE),
				to_sfixed(0.9448,1,L_SIZE),
				to_sfixed(0.9449,1,L_SIZE),
				to_sfixed(0.9449,1,L_SIZE),
				to_sfixed(0.9449,1,L_SIZE),
				to_sfixed(0.9450,1,L_SIZE),
				to_sfixed(0.9450,1,L_SIZE),
				to_sfixed(0.9451,1,L_SIZE),
				to_sfixed(0.9451,1,L_SIZE),
				to_sfixed(0.9451,1,L_SIZE),
				to_sfixed(0.9452,1,L_SIZE),
				to_sfixed(0.9452,1,L_SIZE),
				to_sfixed(0.9453,1,L_SIZE),
				to_sfixed(0.9453,1,L_SIZE),
				to_sfixed(0.9453,1,L_SIZE),
				to_sfixed(0.9454,1,L_SIZE),
				to_sfixed(0.9454,1,L_SIZE),
				to_sfixed(0.9455,1,L_SIZE),
				to_sfixed(0.9455,1,L_SIZE),
				to_sfixed(0.9455,1,L_SIZE),
				to_sfixed(0.9456,1,L_SIZE),
				to_sfixed(0.9456,1,L_SIZE),
				to_sfixed(0.9456,1,L_SIZE),
				to_sfixed(0.9457,1,L_SIZE),
				to_sfixed(0.9457,1,L_SIZE),
				to_sfixed(0.9458,1,L_SIZE),
				to_sfixed(0.9458,1,L_SIZE),
				to_sfixed(0.9458,1,L_SIZE),
				to_sfixed(0.9459,1,L_SIZE),
				to_sfixed(0.9459,1,L_SIZE),
				to_sfixed(0.9460,1,L_SIZE),
				to_sfixed(0.9460,1,L_SIZE),
				to_sfixed(0.9460,1,L_SIZE),
				to_sfixed(0.9461,1,L_SIZE),
				to_sfixed(0.9461,1,L_SIZE),
				to_sfixed(0.9461,1,L_SIZE),
				to_sfixed(0.9462,1,L_SIZE),
				to_sfixed(0.9462,1,L_SIZE),
				to_sfixed(0.9463,1,L_SIZE),
				to_sfixed(0.9463,1,L_SIZE),
				to_sfixed(0.9463,1,L_SIZE),
				to_sfixed(0.9464,1,L_SIZE),
				to_sfixed(0.9464,1,L_SIZE),
				to_sfixed(0.9465,1,L_SIZE),
				to_sfixed(0.9465,1,L_SIZE),
				to_sfixed(0.9465,1,L_SIZE),
				to_sfixed(0.9466,1,L_SIZE),
				to_sfixed(0.9466,1,L_SIZE),
				to_sfixed(0.9466,1,L_SIZE),
				to_sfixed(0.9467,1,L_SIZE),
				to_sfixed(0.9467,1,L_SIZE),
				to_sfixed(0.9468,1,L_SIZE),
				to_sfixed(0.9468,1,L_SIZE),
				to_sfixed(0.9468,1,L_SIZE),
				to_sfixed(0.9469,1,L_SIZE),
				to_sfixed(0.9469,1,L_SIZE),
				to_sfixed(0.9469,1,L_SIZE),
				to_sfixed(0.9470,1,L_SIZE),
				to_sfixed(0.9470,1,L_SIZE),
				to_sfixed(0.9471,1,L_SIZE),
				to_sfixed(0.9471,1,L_SIZE),
				to_sfixed(0.9471,1,L_SIZE),
				to_sfixed(0.9472,1,L_SIZE),
				to_sfixed(0.9472,1,L_SIZE),
				to_sfixed(0.9473,1,L_SIZE),
				to_sfixed(0.9473,1,L_SIZE),
				to_sfixed(0.9473,1,L_SIZE),
				to_sfixed(0.9474,1,L_SIZE),
				to_sfixed(0.9474,1,L_SIZE),
				to_sfixed(0.9474,1,L_SIZE),
				to_sfixed(0.9475,1,L_SIZE),
				to_sfixed(0.9475,1,L_SIZE),
				to_sfixed(0.9476,1,L_SIZE),
				to_sfixed(0.9476,1,L_SIZE),
				to_sfixed(0.9476,1,L_SIZE),
				to_sfixed(0.9477,1,L_SIZE),
				to_sfixed(0.9477,1,L_SIZE),
				to_sfixed(0.9477,1,L_SIZE),
				to_sfixed(0.9478,1,L_SIZE),
				to_sfixed(0.9478,1,L_SIZE),
				to_sfixed(0.9479,1,L_SIZE),
				to_sfixed(0.9479,1,L_SIZE),
				to_sfixed(0.9479,1,L_SIZE),
				to_sfixed(0.9480,1,L_SIZE),
				to_sfixed(0.9480,1,L_SIZE),
				to_sfixed(0.9480,1,L_SIZE),
				to_sfixed(0.9481,1,L_SIZE),
				to_sfixed(0.9481,1,L_SIZE),
				to_sfixed(0.9481,1,L_SIZE),
				to_sfixed(0.9482,1,L_SIZE),
				to_sfixed(0.9482,1,L_SIZE),
				to_sfixed(0.9483,1,L_SIZE),
				to_sfixed(0.9483,1,L_SIZE),
				to_sfixed(0.9483,1,L_SIZE),
				to_sfixed(0.9484,1,L_SIZE),
				to_sfixed(0.9484,1,L_SIZE),
				to_sfixed(0.9484,1,L_SIZE),
				to_sfixed(0.9485,1,L_SIZE),
				to_sfixed(0.9485,1,L_SIZE),
				to_sfixed(0.9486,1,L_SIZE),
				to_sfixed(0.9486,1,L_SIZE),
				to_sfixed(0.9486,1,L_SIZE),
				to_sfixed(0.9487,1,L_SIZE),
				to_sfixed(0.9487,1,L_SIZE),
				to_sfixed(0.9487,1,L_SIZE),
				to_sfixed(0.9488,1,L_SIZE),
				to_sfixed(0.9488,1,L_SIZE),
				to_sfixed(0.9488,1,L_SIZE),
				to_sfixed(0.9489,1,L_SIZE),
				to_sfixed(0.9489,1,L_SIZE),
				to_sfixed(0.9490,1,L_SIZE),
				to_sfixed(0.9490,1,L_SIZE),
				to_sfixed(0.9490,1,L_SIZE),
				to_sfixed(0.9491,1,L_SIZE),
				to_sfixed(0.9491,1,L_SIZE),
				to_sfixed(0.9491,1,L_SIZE),
				to_sfixed(0.9492,1,L_SIZE),
				to_sfixed(0.9492,1,L_SIZE),
				to_sfixed(0.9492,1,L_SIZE),
				to_sfixed(0.9493,1,L_SIZE),
				to_sfixed(0.9493,1,L_SIZE),
				to_sfixed(0.9494,1,L_SIZE),
				to_sfixed(0.9494,1,L_SIZE),
				to_sfixed(0.9494,1,L_SIZE),
				to_sfixed(0.9495,1,L_SIZE),
				to_sfixed(0.9495,1,L_SIZE),
				to_sfixed(0.9495,1,L_SIZE),
				to_sfixed(0.9496,1,L_SIZE),
				to_sfixed(0.9496,1,L_SIZE),
				to_sfixed(0.9496,1,L_SIZE),
				to_sfixed(0.9497,1,L_SIZE),
				to_sfixed(0.9497,1,L_SIZE),
				to_sfixed(0.9498,1,L_SIZE),
				to_sfixed(0.9498,1,L_SIZE),
				to_sfixed(0.9498,1,L_SIZE),
				to_sfixed(0.9499,1,L_SIZE),
				to_sfixed(0.9499,1,L_SIZE),
				to_sfixed(0.9499,1,L_SIZE),
				to_sfixed(0.9500,1,L_SIZE),
				to_sfixed(0.9500,1,L_SIZE),
				to_sfixed(0.9500,1,L_SIZE),
				to_sfixed(0.9501,1,L_SIZE),
				to_sfixed(0.9501,1,L_SIZE),
				to_sfixed(0.9501,1,L_SIZE),
				to_sfixed(0.9502,1,L_SIZE),
				to_sfixed(0.9502,1,L_SIZE),
				to_sfixed(0.9502,1,L_SIZE),
				to_sfixed(0.9503,1,L_SIZE),
				to_sfixed(0.9503,1,L_SIZE),
				to_sfixed(0.9504,1,L_SIZE),
				to_sfixed(0.9504,1,L_SIZE),
				to_sfixed(0.9504,1,L_SIZE),
				to_sfixed(0.9505,1,L_SIZE),
				to_sfixed(0.9505,1,L_SIZE),
				to_sfixed(0.9505,1,L_SIZE),
				to_sfixed(0.9506,1,L_SIZE),
				to_sfixed(0.9506,1,L_SIZE),
				to_sfixed(0.9506,1,L_SIZE),
				to_sfixed(0.9507,1,L_SIZE),
				to_sfixed(0.9507,1,L_SIZE),
				to_sfixed(0.9507,1,L_SIZE),
				to_sfixed(0.9508,1,L_SIZE),
				to_sfixed(0.9508,1,L_SIZE),
				to_sfixed(0.9509,1,L_SIZE),
				to_sfixed(0.9509,1,L_SIZE),
				to_sfixed(0.9509,1,L_SIZE),
				to_sfixed(0.9510,1,L_SIZE),
				to_sfixed(0.9510,1,L_SIZE),
				to_sfixed(0.9510,1,L_SIZE),
				to_sfixed(0.9511,1,L_SIZE),
				to_sfixed(0.9511,1,L_SIZE),
				to_sfixed(0.9511,1,L_SIZE),
				to_sfixed(0.9512,1,L_SIZE),
				to_sfixed(0.9512,1,L_SIZE),
				to_sfixed(0.9512,1,L_SIZE),
				to_sfixed(0.9513,1,L_SIZE),
				to_sfixed(0.9513,1,L_SIZE),
				to_sfixed(0.9513,1,L_SIZE),
				to_sfixed(0.9514,1,L_SIZE),
				to_sfixed(0.9514,1,L_SIZE),
				to_sfixed(0.9514,1,L_SIZE),
				to_sfixed(0.9515,1,L_SIZE),
				to_sfixed(0.9515,1,L_SIZE),
				to_sfixed(0.9515,1,L_SIZE),
				to_sfixed(0.9516,1,L_SIZE),
				to_sfixed(0.9516,1,L_SIZE),
				to_sfixed(0.9517,1,L_SIZE),
				to_sfixed(0.9517,1,L_SIZE),
				to_sfixed(0.9517,1,L_SIZE),
				to_sfixed(0.9518,1,L_SIZE),
				to_sfixed(0.9518,1,L_SIZE),
				to_sfixed(0.9518,1,L_SIZE),
				to_sfixed(0.9519,1,L_SIZE),
				to_sfixed(0.9519,1,L_SIZE),
				to_sfixed(0.9519,1,L_SIZE),
				to_sfixed(0.9520,1,L_SIZE),
				to_sfixed(0.9520,1,L_SIZE),
				to_sfixed(0.9520,1,L_SIZE),
				to_sfixed(0.9521,1,L_SIZE),
				to_sfixed(0.9521,1,L_SIZE),
				to_sfixed(0.9521,1,L_SIZE),
				to_sfixed(0.9522,1,L_SIZE),
				to_sfixed(0.9522,1,L_SIZE),
				to_sfixed(0.9522,1,L_SIZE),
				to_sfixed(0.9523,1,L_SIZE),
				to_sfixed(0.9523,1,L_SIZE),
				to_sfixed(0.9523,1,L_SIZE),
				to_sfixed(0.9524,1,L_SIZE),
				to_sfixed(0.9524,1,L_SIZE),
				to_sfixed(0.9524,1,L_SIZE),
				to_sfixed(0.9525,1,L_SIZE),
				to_sfixed(0.9525,1,L_SIZE),
				to_sfixed(0.9525,1,L_SIZE),
				to_sfixed(0.9526,1,L_SIZE),
				to_sfixed(0.9526,1,L_SIZE),
				to_sfixed(0.9526,1,L_SIZE),
				to_sfixed(0.9527,1,L_SIZE),
				to_sfixed(0.9527,1,L_SIZE),
				to_sfixed(0.9527,1,L_SIZE),
				to_sfixed(0.9528,1,L_SIZE),
				to_sfixed(0.9528,1,L_SIZE),
				to_sfixed(0.9528,1,L_SIZE),
				to_sfixed(0.9529,1,L_SIZE),
				to_sfixed(0.9529,1,L_SIZE),
				to_sfixed(0.9529,1,L_SIZE),
				to_sfixed(0.9530,1,L_SIZE),
				to_sfixed(0.9530,1,L_SIZE),
				to_sfixed(0.9530,1,L_SIZE),
				to_sfixed(0.9531,1,L_SIZE),
				to_sfixed(0.9531,1,L_SIZE),
				to_sfixed(0.9531,1,L_SIZE),
				to_sfixed(0.9532,1,L_SIZE),
				to_sfixed(0.9532,1,L_SIZE),
				to_sfixed(0.9532,1,L_SIZE),
				to_sfixed(0.9533,1,L_SIZE),
				to_sfixed(0.9533,1,L_SIZE),
				to_sfixed(0.9533,1,L_SIZE),
				to_sfixed(0.9534,1,L_SIZE),
				to_sfixed(0.9534,1,L_SIZE),
				to_sfixed(0.9534,1,L_SIZE),
				to_sfixed(0.9535,1,L_SIZE),
				to_sfixed(0.9535,1,L_SIZE),
				to_sfixed(0.9535,1,L_SIZE),
				to_sfixed(0.9536,1,L_SIZE),
				to_sfixed(0.9536,1,L_SIZE),
				to_sfixed(0.9536,1,L_SIZE),
				to_sfixed(0.9537,1,L_SIZE),
				to_sfixed(0.9537,1,L_SIZE),
				to_sfixed(0.9537,1,L_SIZE),
				to_sfixed(0.9538,1,L_SIZE),
				to_sfixed(0.9538,1,L_SIZE),
				to_sfixed(0.9538,1,L_SIZE),
				to_sfixed(0.9539,1,L_SIZE),
				to_sfixed(0.9539,1,L_SIZE),
				to_sfixed(0.9539,1,L_SIZE),
				to_sfixed(0.9540,1,L_SIZE),
				to_sfixed(0.9540,1,L_SIZE),
				to_sfixed(0.9540,1,L_SIZE),
				to_sfixed(0.9541,1,L_SIZE),
				to_sfixed(0.9541,1,L_SIZE),
				to_sfixed(0.9541,1,L_SIZE),
				to_sfixed(0.9542,1,L_SIZE),
				to_sfixed(0.9542,1,L_SIZE),
				to_sfixed(0.9542,1,L_SIZE),
				to_sfixed(0.9543,1,L_SIZE),
				to_sfixed(0.9543,1,L_SIZE),
				to_sfixed(0.9543,1,L_SIZE),
				to_sfixed(0.9544,1,L_SIZE),
				to_sfixed(0.9544,1,L_SIZE),
				to_sfixed(0.9544,1,L_SIZE),
				to_sfixed(0.9545,1,L_SIZE),
				to_sfixed(0.9545,1,L_SIZE),
				to_sfixed(0.9545,1,L_SIZE),
				to_sfixed(0.9546,1,L_SIZE),
				to_sfixed(0.9546,1,L_SIZE),
				to_sfixed(0.9546,1,L_SIZE),
				to_sfixed(0.9547,1,L_SIZE),
				to_sfixed(0.9547,1,L_SIZE),
				to_sfixed(0.9547,1,L_SIZE),
				to_sfixed(0.9548,1,L_SIZE),
				to_sfixed(0.9548,1,L_SIZE),
				to_sfixed(0.9548,1,L_SIZE),
				to_sfixed(0.9549,1,L_SIZE),
				to_sfixed(0.9549,1,L_SIZE),
				to_sfixed(0.9549,1,L_SIZE),
				to_sfixed(0.9550,1,L_SIZE),
				to_sfixed(0.9550,1,L_SIZE),
				to_sfixed(0.9550,1,L_SIZE),
				to_sfixed(0.9551,1,L_SIZE),
				to_sfixed(0.9551,1,L_SIZE),
				to_sfixed(0.9551,1,L_SIZE),
				to_sfixed(0.9552,1,L_SIZE),
				to_sfixed(0.9552,1,L_SIZE),
				to_sfixed(0.9552,1,L_SIZE),
				to_sfixed(0.9552,1,L_SIZE),
				to_sfixed(0.9553,1,L_SIZE),
				to_sfixed(0.9553,1,L_SIZE),
				to_sfixed(0.9553,1,L_SIZE),
				to_sfixed(0.9554,1,L_SIZE),
				to_sfixed(0.9554,1,L_SIZE),
				to_sfixed(0.9554,1,L_SIZE),
				to_sfixed(0.9555,1,L_SIZE),
				to_sfixed(0.9555,1,L_SIZE),
				to_sfixed(0.9555,1,L_SIZE),
				to_sfixed(0.9556,1,L_SIZE),
				to_sfixed(0.9556,1,L_SIZE),
				to_sfixed(0.9556,1,L_SIZE),
				to_sfixed(0.9557,1,L_SIZE),
				to_sfixed(0.9557,1,L_SIZE),
				to_sfixed(0.9557,1,L_SIZE),
				to_sfixed(0.9558,1,L_SIZE),
				to_sfixed(0.9558,1,L_SIZE),
				to_sfixed(0.9558,1,L_SIZE),
				to_sfixed(0.9559,1,L_SIZE),
				to_sfixed(0.9559,1,L_SIZE),
				to_sfixed(0.9559,1,L_SIZE),
				to_sfixed(0.9559,1,L_SIZE),
				to_sfixed(0.9560,1,L_SIZE),
				to_sfixed(0.9560,1,L_SIZE),
				to_sfixed(0.9560,1,L_SIZE),
				to_sfixed(0.9561,1,L_SIZE),
				to_sfixed(0.9561,1,L_SIZE),
				to_sfixed(0.9561,1,L_SIZE),
				to_sfixed(0.9562,1,L_SIZE),
				to_sfixed(0.9562,1,L_SIZE),
				to_sfixed(0.9562,1,L_SIZE),
				to_sfixed(0.9563,1,L_SIZE),
				to_sfixed(0.9563,1,L_SIZE),
				to_sfixed(0.9563,1,L_SIZE),
				to_sfixed(0.9564,1,L_SIZE),
				to_sfixed(0.9564,1,L_SIZE),
				to_sfixed(0.9564,1,L_SIZE),
				to_sfixed(0.9564,1,L_SIZE),
				to_sfixed(0.9565,1,L_SIZE),
				to_sfixed(0.9565,1,L_SIZE),
				to_sfixed(0.9565,1,L_SIZE),
				to_sfixed(0.9566,1,L_SIZE),
				to_sfixed(0.9566,1,L_SIZE),
				to_sfixed(0.9566,1,L_SIZE),
				to_sfixed(0.9567,1,L_SIZE),
				to_sfixed(0.9567,1,L_SIZE),
				to_sfixed(0.9567,1,L_SIZE),
				to_sfixed(0.9568,1,L_SIZE),
				to_sfixed(0.9568,1,L_SIZE),
				to_sfixed(0.9568,1,L_SIZE),
				to_sfixed(0.9569,1,L_SIZE),
				to_sfixed(0.9569,1,L_SIZE),
				to_sfixed(0.9569,1,L_SIZE),
				to_sfixed(0.9569,1,L_SIZE),
				to_sfixed(0.9570,1,L_SIZE),
				to_sfixed(0.9570,1,L_SIZE),
				to_sfixed(0.9570,1,L_SIZE),
				to_sfixed(0.9571,1,L_SIZE),
				to_sfixed(0.9571,1,L_SIZE),
				to_sfixed(0.9571,1,L_SIZE),
				to_sfixed(0.9572,1,L_SIZE),
				to_sfixed(0.9572,1,L_SIZE),
				to_sfixed(0.9572,1,L_SIZE),
				to_sfixed(0.9573,1,L_SIZE),
				to_sfixed(0.9573,1,L_SIZE),
				to_sfixed(0.9573,1,L_SIZE),
				to_sfixed(0.9573,1,L_SIZE),
				to_sfixed(0.9574,1,L_SIZE),
				to_sfixed(0.9574,1,L_SIZE),
				to_sfixed(0.9574,1,L_SIZE),
				to_sfixed(0.9575,1,L_SIZE),
				to_sfixed(0.9575,1,L_SIZE),
				to_sfixed(0.9575,1,L_SIZE),
				to_sfixed(0.9576,1,L_SIZE),
				to_sfixed(0.9576,1,L_SIZE),
				to_sfixed(0.9576,1,L_SIZE),
				to_sfixed(0.9576,1,L_SIZE),
				to_sfixed(0.9577,1,L_SIZE),
				to_sfixed(0.9577,1,L_SIZE),
				to_sfixed(0.9577,1,L_SIZE),
				to_sfixed(0.9578,1,L_SIZE),
				to_sfixed(0.9578,1,L_SIZE),
				to_sfixed(0.9578,1,L_SIZE),
				to_sfixed(0.9579,1,L_SIZE),
				to_sfixed(0.9579,1,L_SIZE),
				to_sfixed(0.9579,1,L_SIZE),
				to_sfixed(0.9580,1,L_SIZE),
				to_sfixed(0.9580,1,L_SIZE),
				to_sfixed(0.9580,1,L_SIZE),
				to_sfixed(0.9580,1,L_SIZE),
				to_sfixed(0.9581,1,L_SIZE),
				to_sfixed(0.9581,1,L_SIZE),
				to_sfixed(0.9581,1,L_SIZE),
				to_sfixed(0.9582,1,L_SIZE),
				to_sfixed(0.9582,1,L_SIZE),
				to_sfixed(0.9582,1,L_SIZE),
				to_sfixed(0.9583,1,L_SIZE),
				to_sfixed(0.9583,1,L_SIZE),
				to_sfixed(0.9583,1,L_SIZE),
				to_sfixed(0.9583,1,L_SIZE),
				to_sfixed(0.9584,1,L_SIZE),
				to_sfixed(0.9584,1,L_SIZE),
				to_sfixed(0.9584,1,L_SIZE),
				to_sfixed(0.9585,1,L_SIZE),
				to_sfixed(0.9585,1,L_SIZE),
				to_sfixed(0.9585,1,L_SIZE),
				to_sfixed(0.9585,1,L_SIZE),
				to_sfixed(0.9586,1,L_SIZE),
				to_sfixed(0.9586,1,L_SIZE),
				to_sfixed(0.9586,1,L_SIZE),
				to_sfixed(0.9587,1,L_SIZE),
				to_sfixed(0.9587,1,L_SIZE),
				to_sfixed(0.9587,1,L_SIZE),
				to_sfixed(0.9588,1,L_SIZE),
				to_sfixed(0.9588,1,L_SIZE),
				to_sfixed(0.9588,1,L_SIZE),
				to_sfixed(0.9588,1,L_SIZE),
				to_sfixed(0.9589,1,L_SIZE),
				to_sfixed(0.9589,1,L_SIZE),
				to_sfixed(0.9589,1,L_SIZE),
				to_sfixed(0.9590,1,L_SIZE),
				to_sfixed(0.9590,1,L_SIZE),
				to_sfixed(0.9590,1,L_SIZE),
				to_sfixed(0.9591,1,L_SIZE),
				to_sfixed(0.9591,1,L_SIZE),
				to_sfixed(0.9591,1,L_SIZE),
				to_sfixed(0.9591,1,L_SIZE),
				to_sfixed(0.9592,1,L_SIZE),
				to_sfixed(0.9592,1,L_SIZE),
				to_sfixed(0.9592,1,L_SIZE),
				to_sfixed(0.9593,1,L_SIZE),
				to_sfixed(0.9593,1,L_SIZE),
				to_sfixed(0.9593,1,L_SIZE),
				to_sfixed(0.9593,1,L_SIZE),
				to_sfixed(0.9594,1,L_SIZE),
				to_sfixed(0.9594,1,L_SIZE),
				to_sfixed(0.9594,1,L_SIZE),
				to_sfixed(0.9595,1,L_SIZE),
				to_sfixed(0.9595,1,L_SIZE),
				to_sfixed(0.9595,1,L_SIZE),
				to_sfixed(0.9595,1,L_SIZE),
				to_sfixed(0.9596,1,L_SIZE),
				to_sfixed(0.9596,1,L_SIZE),
				to_sfixed(0.9596,1,L_SIZE),
				to_sfixed(0.9597,1,L_SIZE),
				to_sfixed(0.9597,1,L_SIZE),
				to_sfixed(0.9597,1,L_SIZE),
				to_sfixed(0.9598,1,L_SIZE),
				to_sfixed(0.9598,1,L_SIZE),
				to_sfixed(0.9598,1,L_SIZE),
				to_sfixed(0.9598,1,L_SIZE),
				to_sfixed(0.9599,1,L_SIZE),
				to_sfixed(0.9599,1,L_SIZE),
				to_sfixed(0.9599,1,L_SIZE),
				to_sfixed(0.9600,1,L_SIZE),
				to_sfixed(0.9600,1,L_SIZE),
				to_sfixed(0.9600,1,L_SIZE),
				to_sfixed(0.9600,1,L_SIZE),
				to_sfixed(0.9601,1,L_SIZE),
				to_sfixed(0.9601,1,L_SIZE),
				to_sfixed(0.9601,1,L_SIZE),
				to_sfixed(0.9602,1,L_SIZE),
				to_sfixed(0.9602,1,L_SIZE),
				to_sfixed(0.9602,1,L_SIZE),
				to_sfixed(0.9602,1,L_SIZE),
				to_sfixed(0.9603,1,L_SIZE),
				to_sfixed(0.9603,1,L_SIZE),
				to_sfixed(0.9603,1,L_SIZE),
				to_sfixed(0.9604,1,L_SIZE),
				to_sfixed(0.9604,1,L_SIZE),
				to_sfixed(0.9604,1,L_SIZE),
				to_sfixed(0.9604,1,L_SIZE),
				to_sfixed(0.9605,1,L_SIZE),
				to_sfixed(0.9605,1,L_SIZE),
				to_sfixed(0.9605,1,L_SIZE),
				to_sfixed(0.9606,1,L_SIZE),
				to_sfixed(0.9606,1,L_SIZE),
				to_sfixed(0.9606,1,L_SIZE),
				to_sfixed(0.9606,1,L_SIZE),
				to_sfixed(0.9607,1,L_SIZE),
				to_sfixed(0.9607,1,L_SIZE),
				to_sfixed(0.9607,1,L_SIZE),
				to_sfixed(0.9608,1,L_SIZE),
				to_sfixed(0.9608,1,L_SIZE),
				to_sfixed(0.9608,1,L_SIZE),
				to_sfixed(0.9608,1,L_SIZE),
				to_sfixed(0.9609,1,L_SIZE),
				to_sfixed(0.9609,1,L_SIZE),
				to_sfixed(0.9609,1,L_SIZE),
				to_sfixed(0.9609,1,L_SIZE),
				to_sfixed(0.9610,1,L_SIZE),
				to_sfixed(0.9610,1,L_SIZE),
				to_sfixed(0.9610,1,L_SIZE),
				to_sfixed(0.9611,1,L_SIZE),
				to_sfixed(0.9611,1,L_SIZE),
				to_sfixed(0.9611,1,L_SIZE),
				to_sfixed(0.9611,1,L_SIZE),
				to_sfixed(0.9612,1,L_SIZE),
				to_sfixed(0.9612,1,L_SIZE),
				to_sfixed(0.9612,1,L_SIZE),
				to_sfixed(0.9613,1,L_SIZE),
				to_sfixed(0.9613,1,L_SIZE),
				to_sfixed(0.9613,1,L_SIZE),
				to_sfixed(0.9613,1,L_SIZE),
				to_sfixed(0.9614,1,L_SIZE),
				to_sfixed(0.9614,1,L_SIZE),
				to_sfixed(0.9614,1,L_SIZE),
				to_sfixed(0.9614,1,L_SIZE),
				to_sfixed(0.9615,1,L_SIZE),
				to_sfixed(0.9615,1,L_SIZE),
				to_sfixed(0.9615,1,L_SIZE),
				to_sfixed(0.9616,1,L_SIZE),
				to_sfixed(0.9616,1,L_SIZE),
				to_sfixed(0.9616,1,L_SIZE),
				to_sfixed(0.9616,1,L_SIZE),
				to_sfixed(0.9617,1,L_SIZE),
				to_sfixed(0.9617,1,L_SIZE),
				to_sfixed(0.9617,1,L_SIZE),
				to_sfixed(0.9618,1,L_SIZE),
				to_sfixed(0.9618,1,L_SIZE),
				to_sfixed(0.9618,1,L_SIZE),
				to_sfixed(0.9618,1,L_SIZE),
				to_sfixed(0.9619,1,L_SIZE),
				to_sfixed(0.9619,1,L_SIZE),
				to_sfixed(0.9619,1,L_SIZE),
				to_sfixed(0.9619,1,L_SIZE),
				to_sfixed(0.9620,1,L_SIZE),
				to_sfixed(0.9620,1,L_SIZE),
				to_sfixed(0.9620,1,L_SIZE),
				to_sfixed(0.9621,1,L_SIZE),
				to_sfixed(0.9621,1,L_SIZE),
				to_sfixed(0.9621,1,L_SIZE),
				to_sfixed(0.9621,1,L_SIZE),
				to_sfixed(0.9622,1,L_SIZE),
				to_sfixed(0.9622,1,L_SIZE),
				to_sfixed(0.9622,1,L_SIZE),
				to_sfixed(0.9622,1,L_SIZE),
				to_sfixed(0.9623,1,L_SIZE),
				to_sfixed(0.9623,1,L_SIZE),
				to_sfixed(0.9623,1,L_SIZE),
				to_sfixed(0.9624,1,L_SIZE),
				to_sfixed(0.9624,1,L_SIZE),
				to_sfixed(0.9624,1,L_SIZE),
				to_sfixed(0.9624,1,L_SIZE),
				to_sfixed(0.9625,1,L_SIZE),
				to_sfixed(0.9625,1,L_SIZE),
				to_sfixed(0.9625,1,L_SIZE),
				to_sfixed(0.9625,1,L_SIZE),
				to_sfixed(0.9626,1,L_SIZE),
				to_sfixed(0.9626,1,L_SIZE),
				to_sfixed(0.9626,1,L_SIZE),
				to_sfixed(0.9626,1,L_SIZE),
				to_sfixed(0.9627,1,L_SIZE),
				to_sfixed(0.9627,1,L_SIZE),
				to_sfixed(0.9627,1,L_SIZE),
				to_sfixed(0.9628,1,L_SIZE),
				to_sfixed(0.9628,1,L_SIZE),
				to_sfixed(0.9628,1,L_SIZE),
				to_sfixed(0.9628,1,L_SIZE),
				to_sfixed(0.9629,1,L_SIZE),
				to_sfixed(0.9629,1,L_SIZE),
				to_sfixed(0.9629,1,L_SIZE),
				to_sfixed(0.9629,1,L_SIZE),
				to_sfixed(0.9630,1,L_SIZE),
				to_sfixed(0.9630,1,L_SIZE),
				to_sfixed(0.9630,1,L_SIZE),
				to_sfixed(0.9630,1,L_SIZE),
				to_sfixed(0.9631,1,L_SIZE),
				to_sfixed(0.9631,1,L_SIZE),
				to_sfixed(0.9631,1,L_SIZE),
				to_sfixed(0.9632,1,L_SIZE),
				to_sfixed(0.9632,1,L_SIZE),
				to_sfixed(0.9632,1,L_SIZE),
				to_sfixed(0.9632,1,L_SIZE),
				to_sfixed(0.9633,1,L_SIZE),
				to_sfixed(0.9633,1,L_SIZE),
				to_sfixed(0.9633,1,L_SIZE),
				to_sfixed(0.9633,1,L_SIZE),
				to_sfixed(0.9634,1,L_SIZE),
				to_sfixed(0.9634,1,L_SIZE),
				to_sfixed(0.9634,1,L_SIZE),
				to_sfixed(0.9634,1,L_SIZE),
				to_sfixed(0.9635,1,L_SIZE),
				to_sfixed(0.9635,1,L_SIZE),
				to_sfixed(0.9635,1,L_SIZE),
				to_sfixed(0.9636,1,L_SIZE),
				to_sfixed(0.9636,1,L_SIZE),
				to_sfixed(0.9636,1,L_SIZE),
				to_sfixed(0.9636,1,L_SIZE),
				to_sfixed(0.9637,1,L_SIZE),
				to_sfixed(0.9637,1,L_SIZE),
				to_sfixed(0.9637,1,L_SIZE),
				to_sfixed(0.9637,1,L_SIZE),
				to_sfixed(0.9638,1,L_SIZE),
				to_sfixed(0.9638,1,L_SIZE),
				to_sfixed(0.9638,1,L_SIZE),
				to_sfixed(0.9638,1,L_SIZE),
				to_sfixed(0.9639,1,L_SIZE),
				to_sfixed(0.9639,1,L_SIZE),
				to_sfixed(0.9639,1,L_SIZE),
				to_sfixed(0.9639,1,L_SIZE),
				to_sfixed(0.9640,1,L_SIZE),
				to_sfixed(0.9640,1,L_SIZE),
				to_sfixed(0.9640,1,L_SIZE),
				to_sfixed(0.9640,1,L_SIZE),
				to_sfixed(0.9641,1,L_SIZE),
				to_sfixed(0.9641,1,L_SIZE),
				to_sfixed(0.9641,1,L_SIZE),
				to_sfixed(0.9641,1,L_SIZE),
				to_sfixed(0.9642,1,L_SIZE),
				to_sfixed(0.9642,1,L_SIZE),
				to_sfixed(0.9642,1,L_SIZE),
				to_sfixed(0.9643,1,L_SIZE),
				to_sfixed(0.9643,1,L_SIZE),
				to_sfixed(0.9643,1,L_SIZE),
				to_sfixed(0.9643,1,L_SIZE),
				to_sfixed(0.9644,1,L_SIZE),
				to_sfixed(0.9644,1,L_SIZE),
				to_sfixed(0.9644,1,L_SIZE),
				to_sfixed(0.9644,1,L_SIZE),
				to_sfixed(0.9645,1,L_SIZE),
				to_sfixed(0.9645,1,L_SIZE),
				to_sfixed(0.9645,1,L_SIZE),
				to_sfixed(0.9645,1,L_SIZE),
				to_sfixed(0.9646,1,L_SIZE),
				to_sfixed(0.9646,1,L_SIZE),
				to_sfixed(0.9646,1,L_SIZE),
				to_sfixed(0.9646,1,L_SIZE),
				to_sfixed(0.9647,1,L_SIZE),
				to_sfixed(0.9647,1,L_SIZE),
				to_sfixed(0.9647,1,L_SIZE),
				to_sfixed(0.9647,1,L_SIZE),
				to_sfixed(0.9648,1,L_SIZE),
				to_sfixed(0.9648,1,L_SIZE),
				to_sfixed(0.9648,1,L_SIZE),
				to_sfixed(0.9648,1,L_SIZE),
				to_sfixed(0.9649,1,L_SIZE),
				to_sfixed(0.9649,1,L_SIZE),
				to_sfixed(0.9649,1,L_SIZE),
				to_sfixed(0.9649,1,L_SIZE),
				to_sfixed(0.9650,1,L_SIZE),
				to_sfixed(0.9650,1,L_SIZE),
				to_sfixed(0.9650,1,L_SIZE),
				to_sfixed(0.9650,1,L_SIZE),
				to_sfixed(0.9651,1,L_SIZE),
				to_sfixed(0.9651,1,L_SIZE),
				to_sfixed(0.9651,1,L_SIZE),
				to_sfixed(0.9651,1,L_SIZE),
				to_sfixed(0.9652,1,L_SIZE),
				to_sfixed(0.9652,1,L_SIZE),
				to_sfixed(0.9652,1,L_SIZE),
				to_sfixed(0.9652,1,L_SIZE),
				to_sfixed(0.9653,1,L_SIZE),
				to_sfixed(0.9653,1,L_SIZE),
				to_sfixed(0.9653,1,L_SIZE),
				to_sfixed(0.9653,1,L_SIZE),
				to_sfixed(0.9654,1,L_SIZE),
				to_sfixed(0.9654,1,L_SIZE),
				to_sfixed(0.9654,1,L_SIZE),
				to_sfixed(0.9654,1,L_SIZE),
				to_sfixed(0.9655,1,L_SIZE),
				to_sfixed(0.9655,1,L_SIZE),
				to_sfixed(0.9655,1,L_SIZE),
				to_sfixed(0.9655,1,L_SIZE),
				to_sfixed(0.9656,1,L_SIZE),
				to_sfixed(0.9656,1,L_SIZE),
				to_sfixed(0.9656,1,L_SIZE),
				to_sfixed(0.9656,1,L_SIZE),
				to_sfixed(0.9657,1,L_SIZE),
				to_sfixed(0.9657,1,L_SIZE),
				to_sfixed(0.9657,1,L_SIZE),
				to_sfixed(0.9657,1,L_SIZE),
				to_sfixed(0.9658,1,L_SIZE),
				to_sfixed(0.9658,1,L_SIZE),
				to_sfixed(0.9658,1,L_SIZE),
				to_sfixed(0.9658,1,L_SIZE),
				to_sfixed(0.9659,1,L_SIZE),
				to_sfixed(0.9659,1,L_SIZE),
				to_sfixed(0.9659,1,L_SIZE),
				to_sfixed(0.9659,1,L_SIZE),
				to_sfixed(0.9660,1,L_SIZE),
				to_sfixed(0.9660,1,L_SIZE),
				to_sfixed(0.9660,1,L_SIZE),
				to_sfixed(0.9660,1,L_SIZE),
				to_sfixed(0.9661,1,L_SIZE),
				to_sfixed(0.9661,1,L_SIZE),
				to_sfixed(0.9661,1,L_SIZE),
				to_sfixed(0.9661,1,L_SIZE),
				to_sfixed(0.9662,1,L_SIZE),
				to_sfixed(0.9662,1,L_SIZE),
				to_sfixed(0.9662,1,L_SIZE),
				to_sfixed(0.9662,1,L_SIZE),
				to_sfixed(0.9663,1,L_SIZE),
				to_sfixed(0.9663,1,L_SIZE),
				to_sfixed(0.9663,1,L_SIZE),
				to_sfixed(0.9663,1,L_SIZE),
				to_sfixed(0.9663,1,L_SIZE),
				to_sfixed(0.9664,1,L_SIZE),
				to_sfixed(0.9664,1,L_SIZE),
				to_sfixed(0.9664,1,L_SIZE),
				to_sfixed(0.9664,1,L_SIZE),
				to_sfixed(0.9665,1,L_SIZE),
				to_sfixed(0.9665,1,L_SIZE),
				to_sfixed(0.9665,1,L_SIZE),
				to_sfixed(0.9665,1,L_SIZE),
				to_sfixed(0.9666,1,L_SIZE),
				to_sfixed(0.9666,1,L_SIZE),
				to_sfixed(0.9666,1,L_SIZE),
				to_sfixed(0.9666,1,L_SIZE),
				to_sfixed(0.9667,1,L_SIZE),
				to_sfixed(0.9667,1,L_SIZE),
				to_sfixed(0.9667,1,L_SIZE),
				to_sfixed(0.9667,1,L_SIZE),
				to_sfixed(0.9668,1,L_SIZE),
				to_sfixed(0.9668,1,L_SIZE),
				to_sfixed(0.9668,1,L_SIZE),
				to_sfixed(0.9668,1,L_SIZE),
				to_sfixed(0.9669,1,L_SIZE),
				to_sfixed(0.9669,1,L_SIZE),
				to_sfixed(0.9669,1,L_SIZE),
				to_sfixed(0.9669,1,L_SIZE),
				to_sfixed(0.9669,1,L_SIZE),
				to_sfixed(0.9670,1,L_SIZE),
				to_sfixed(0.9670,1,L_SIZE),
				to_sfixed(0.9670,1,L_SIZE),
				to_sfixed(0.9670,1,L_SIZE),
				to_sfixed(0.9671,1,L_SIZE),
				to_sfixed(0.9671,1,L_SIZE),
				to_sfixed(0.9671,1,L_SIZE),
				to_sfixed(0.9671,1,L_SIZE),
				to_sfixed(0.9672,1,L_SIZE),
				to_sfixed(0.9672,1,L_SIZE),
				to_sfixed(0.9672,1,L_SIZE),
				to_sfixed(0.9672,1,L_SIZE),
				to_sfixed(0.9673,1,L_SIZE),
				to_sfixed(0.9673,1,L_SIZE),
				to_sfixed(0.9673,1,L_SIZE),
				to_sfixed(0.9673,1,L_SIZE),
				to_sfixed(0.9674,1,L_SIZE),
				to_sfixed(0.9674,1,L_SIZE),
				to_sfixed(0.9674,1,L_SIZE),
				to_sfixed(0.9674,1,L_SIZE),
				to_sfixed(0.9674,1,L_SIZE),
				to_sfixed(0.9675,1,L_SIZE),
				to_sfixed(0.9675,1,L_SIZE),
				to_sfixed(0.9675,1,L_SIZE),
				to_sfixed(0.9675,1,L_SIZE),
				to_sfixed(0.9676,1,L_SIZE),
				to_sfixed(0.9676,1,L_SIZE),
				to_sfixed(0.9676,1,L_SIZE),
				to_sfixed(0.9676,1,L_SIZE),
				to_sfixed(0.9677,1,L_SIZE),
				to_sfixed(0.9677,1,L_SIZE),
				to_sfixed(0.9677,1,L_SIZE),
				to_sfixed(0.9677,1,L_SIZE),
				to_sfixed(0.9677,1,L_SIZE),
				to_sfixed(0.9678,1,L_SIZE),
				to_sfixed(0.9678,1,L_SIZE),
				to_sfixed(0.9678,1,L_SIZE),
				to_sfixed(0.9678,1,L_SIZE),
				to_sfixed(0.9679,1,L_SIZE),
				to_sfixed(0.9679,1,L_SIZE),
				to_sfixed(0.9679,1,L_SIZE),
				to_sfixed(0.9679,1,L_SIZE),
				to_sfixed(0.9680,1,L_SIZE),
				to_sfixed(0.9680,1,L_SIZE),
				to_sfixed(0.9680,1,L_SIZE),
				to_sfixed(0.9680,1,L_SIZE),
				to_sfixed(0.9680,1,L_SIZE),
				to_sfixed(0.9681,1,L_SIZE),
				to_sfixed(0.9681,1,L_SIZE),
				to_sfixed(0.9681,1,L_SIZE),
				to_sfixed(0.9681,1,L_SIZE),
				to_sfixed(0.9682,1,L_SIZE),
				to_sfixed(0.9682,1,L_SIZE),
				to_sfixed(0.9682,1,L_SIZE),
				to_sfixed(0.9682,1,L_SIZE),
				to_sfixed(0.9683,1,L_SIZE),
				to_sfixed(0.9683,1,L_SIZE),
				to_sfixed(0.9683,1,L_SIZE),
				to_sfixed(0.9683,1,L_SIZE),
				to_sfixed(0.9683,1,L_SIZE),
				to_sfixed(0.9684,1,L_SIZE),
				to_sfixed(0.9684,1,L_SIZE),
				to_sfixed(0.9684,1,L_SIZE),
				to_sfixed(0.9684,1,L_SIZE),
				to_sfixed(0.9685,1,L_SIZE),
				to_sfixed(0.9685,1,L_SIZE),
				to_sfixed(0.9685,1,L_SIZE),
				to_sfixed(0.9685,1,L_SIZE),
				to_sfixed(0.9686,1,L_SIZE),
				to_sfixed(0.9686,1,L_SIZE),
				to_sfixed(0.9686,1,L_SIZE),
				to_sfixed(0.9686,1,L_SIZE),
				to_sfixed(0.9686,1,L_SIZE),
				to_sfixed(0.9687,1,L_SIZE),
				to_sfixed(0.9687,1,L_SIZE),
				to_sfixed(0.9687,1,L_SIZE),
				to_sfixed(0.9687,1,L_SIZE),
				to_sfixed(0.9688,1,L_SIZE),
				to_sfixed(0.9688,1,L_SIZE),
				to_sfixed(0.9688,1,L_SIZE),
				to_sfixed(0.9688,1,L_SIZE),
				to_sfixed(0.9688,1,L_SIZE),
				to_sfixed(0.9689,1,L_SIZE),
				to_sfixed(0.9689,1,L_SIZE),
				to_sfixed(0.9689,1,L_SIZE),
				to_sfixed(0.9689,1,L_SIZE),
				to_sfixed(0.9690,1,L_SIZE),
				to_sfixed(0.9690,1,L_SIZE),
				to_sfixed(0.9690,1,L_SIZE),
				to_sfixed(0.9690,1,L_SIZE),
				to_sfixed(0.9690,1,L_SIZE),
				to_sfixed(0.9691,1,L_SIZE),
				to_sfixed(0.9691,1,L_SIZE),
				to_sfixed(0.9691,1,L_SIZE),
				to_sfixed(0.9691,1,L_SIZE),
				to_sfixed(0.9692,1,L_SIZE),
				to_sfixed(0.9692,1,L_SIZE),
				to_sfixed(0.9692,1,L_SIZE),
				to_sfixed(0.9692,1,L_SIZE),
				to_sfixed(0.9692,1,L_SIZE),
				to_sfixed(0.9693,1,L_SIZE),
				to_sfixed(0.9693,1,L_SIZE),
				to_sfixed(0.9693,1,L_SIZE),
				to_sfixed(0.9693,1,L_SIZE),
				to_sfixed(0.9694,1,L_SIZE),
				to_sfixed(0.9694,1,L_SIZE),
				to_sfixed(0.9694,1,L_SIZE),
				to_sfixed(0.9694,1,L_SIZE),
				to_sfixed(0.9694,1,L_SIZE),
				to_sfixed(0.9695,1,L_SIZE),
				to_sfixed(0.9695,1,L_SIZE),
				to_sfixed(0.9695,1,L_SIZE),
				to_sfixed(0.9695,1,L_SIZE),
				to_sfixed(0.9696,1,L_SIZE),
				to_sfixed(0.9696,1,L_SIZE),
				to_sfixed(0.9696,1,L_SIZE),
				to_sfixed(0.9696,1,L_SIZE),
				to_sfixed(0.9696,1,L_SIZE),
				to_sfixed(0.9697,1,L_SIZE),
				to_sfixed(0.9697,1,L_SIZE),
				to_sfixed(0.9697,1,L_SIZE),
				to_sfixed(0.9697,1,L_SIZE),
				to_sfixed(0.9698,1,L_SIZE),
				to_sfixed(0.9698,1,L_SIZE),
				to_sfixed(0.9698,1,L_SIZE),
				to_sfixed(0.9698,1,L_SIZE),
				to_sfixed(0.9698,1,L_SIZE),
				to_sfixed(0.9699,1,L_SIZE),
				to_sfixed(0.9699,1,L_SIZE),
				to_sfixed(0.9699,1,L_SIZE),
				to_sfixed(0.9699,1,L_SIZE),
				to_sfixed(0.9699,1,L_SIZE),
				to_sfixed(0.9700,1,L_SIZE),
				to_sfixed(0.9700,1,L_SIZE),
				to_sfixed(0.9700,1,L_SIZE),
				to_sfixed(0.9700,1,L_SIZE),
				to_sfixed(0.9701,1,L_SIZE),
				to_sfixed(0.9701,1,L_SIZE),
				to_sfixed(0.9701,1,L_SIZE),
				to_sfixed(0.9701,1,L_SIZE),
				to_sfixed(0.9701,1,L_SIZE),
				to_sfixed(0.9702,1,L_SIZE),
				to_sfixed(0.9702,1,L_SIZE),
				to_sfixed(0.9702,1,L_SIZE),
				to_sfixed(0.9702,1,L_SIZE),
				to_sfixed(0.9703,1,L_SIZE),
				to_sfixed(0.9703,1,L_SIZE),
				to_sfixed(0.9703,1,L_SIZE),
				to_sfixed(0.9703,1,L_SIZE),
				to_sfixed(0.9703,1,L_SIZE),
				to_sfixed(0.9704,1,L_SIZE),
				to_sfixed(0.9704,1,L_SIZE),
				to_sfixed(0.9704,1,L_SIZE),
				to_sfixed(0.9704,1,L_SIZE),
				to_sfixed(0.9704,1,L_SIZE),
				to_sfixed(0.9705,1,L_SIZE),
				to_sfixed(0.9705,1,L_SIZE),
				to_sfixed(0.9705,1,L_SIZE),
				to_sfixed(0.9705,1,L_SIZE),
				to_sfixed(0.9705,1,L_SIZE),
				to_sfixed(0.9706,1,L_SIZE),
				to_sfixed(0.9706,1,L_SIZE),
				to_sfixed(0.9706,1,L_SIZE),
				to_sfixed(0.9706,1,L_SIZE),
				to_sfixed(0.9707,1,L_SIZE),
				to_sfixed(0.9707,1,L_SIZE),
				to_sfixed(0.9707,1,L_SIZE),
				to_sfixed(0.9707,1,L_SIZE),
				to_sfixed(0.9707,1,L_SIZE),
				to_sfixed(0.9708,1,L_SIZE),
				to_sfixed(0.9708,1,L_SIZE),
				to_sfixed(0.9708,1,L_SIZE),
				to_sfixed(0.9708,1,L_SIZE),
				to_sfixed(0.9708,1,L_SIZE),
				to_sfixed(0.9709,1,L_SIZE),
				to_sfixed(0.9709,1,L_SIZE),
				to_sfixed(0.9709,1,L_SIZE),
				to_sfixed(0.9709,1,L_SIZE),
				to_sfixed(0.9710,1,L_SIZE),
				to_sfixed(0.9710,1,L_SIZE),
				to_sfixed(0.9710,1,L_SIZE),
				to_sfixed(0.9710,1,L_SIZE),
				to_sfixed(0.9710,1,L_SIZE),
				to_sfixed(0.9711,1,L_SIZE),
				to_sfixed(0.9711,1,L_SIZE),
				to_sfixed(0.9711,1,L_SIZE),
				to_sfixed(0.9711,1,L_SIZE),
				to_sfixed(0.9711,1,L_SIZE),
				to_sfixed(0.9712,1,L_SIZE),
				to_sfixed(0.9712,1,L_SIZE),
				to_sfixed(0.9712,1,L_SIZE),
				to_sfixed(0.9712,1,L_SIZE),
				to_sfixed(0.9712,1,L_SIZE),
				to_sfixed(0.9713,1,L_SIZE),
				to_sfixed(0.9713,1,L_SIZE),
				to_sfixed(0.9713,1,L_SIZE),
				to_sfixed(0.9713,1,L_SIZE),
				to_sfixed(0.9713,1,L_SIZE),
				to_sfixed(0.9714,1,L_SIZE),
				to_sfixed(0.9714,1,L_SIZE),
				to_sfixed(0.9714,1,L_SIZE),
				to_sfixed(0.9714,1,L_SIZE),
				to_sfixed(0.9714,1,L_SIZE),
				to_sfixed(0.9715,1,L_SIZE),
				to_sfixed(0.9715,1,L_SIZE),
				to_sfixed(0.9715,1,L_SIZE),
				to_sfixed(0.9715,1,L_SIZE),
				to_sfixed(0.9716,1,L_SIZE),
				to_sfixed(0.9716,1,L_SIZE),
				to_sfixed(0.9716,1,L_SIZE),
				to_sfixed(0.9716,1,L_SIZE),
				to_sfixed(0.9716,1,L_SIZE),
				to_sfixed(0.9717,1,L_SIZE),
				to_sfixed(0.9717,1,L_SIZE),
				to_sfixed(0.9717,1,L_SIZE),
				to_sfixed(0.9717,1,L_SIZE),
				to_sfixed(0.9717,1,L_SIZE),
				to_sfixed(0.9718,1,L_SIZE),
				to_sfixed(0.9718,1,L_SIZE),
				to_sfixed(0.9718,1,L_SIZE),
				to_sfixed(0.9718,1,L_SIZE),
				to_sfixed(0.9718,1,L_SIZE),
				to_sfixed(0.9719,1,L_SIZE),
				to_sfixed(0.9719,1,L_SIZE),
				to_sfixed(0.9719,1,L_SIZE),
				to_sfixed(0.9719,1,L_SIZE),
				to_sfixed(0.9719,1,L_SIZE),
				to_sfixed(0.9720,1,L_SIZE),
				to_sfixed(0.9720,1,L_SIZE),
				to_sfixed(0.9720,1,L_SIZE),
				to_sfixed(0.9720,1,L_SIZE),
				to_sfixed(0.9720,1,L_SIZE),
				to_sfixed(0.9721,1,L_SIZE),
				to_sfixed(0.9721,1,L_SIZE),
				to_sfixed(0.9721,1,L_SIZE),
				to_sfixed(0.9721,1,L_SIZE),
				to_sfixed(0.9721,1,L_SIZE),
				to_sfixed(0.9722,1,L_SIZE),
				to_sfixed(0.9722,1,L_SIZE),
				to_sfixed(0.9722,1,L_SIZE),
				to_sfixed(0.9722,1,L_SIZE),
				to_sfixed(0.9722,1,L_SIZE),
				to_sfixed(0.9723,1,L_SIZE),
				to_sfixed(0.9723,1,L_SIZE),
				to_sfixed(0.9723,1,L_SIZE),
				to_sfixed(0.9723,1,L_SIZE),
				to_sfixed(0.9723,1,L_SIZE),
				to_sfixed(0.9724,1,L_SIZE),
				to_sfixed(0.9724,1,L_SIZE),
				to_sfixed(0.9724,1,L_SIZE),
				to_sfixed(0.9724,1,L_SIZE),
				to_sfixed(0.9724,1,L_SIZE),
				to_sfixed(0.9725,1,L_SIZE),
				to_sfixed(0.9725,1,L_SIZE),
				to_sfixed(0.9725,1,L_SIZE),
				to_sfixed(0.9725,1,L_SIZE),
				to_sfixed(0.9725,1,L_SIZE),
				to_sfixed(0.9726,1,L_SIZE),
				to_sfixed(0.9726,1,L_SIZE),
				to_sfixed(0.9726,1,L_SIZE),
				to_sfixed(0.9726,1,L_SIZE),
				to_sfixed(0.9726,1,L_SIZE),
				to_sfixed(0.9727,1,L_SIZE),
				to_sfixed(0.9727,1,L_SIZE),
				to_sfixed(0.9727,1,L_SIZE),
				to_sfixed(0.9727,1,L_SIZE),
				to_sfixed(0.9727,1,L_SIZE),
				to_sfixed(0.9728,1,L_SIZE),
				to_sfixed(0.9728,1,L_SIZE),
				to_sfixed(0.9728,1,L_SIZE),
				to_sfixed(0.9728,1,L_SIZE),
				to_sfixed(0.9728,1,L_SIZE),
				to_sfixed(0.9729,1,L_SIZE),
				to_sfixed(0.9729,1,L_SIZE),
				to_sfixed(0.9729,1,L_SIZE),
				to_sfixed(0.9729,1,L_SIZE),
				to_sfixed(0.9729,1,L_SIZE),
				to_sfixed(0.9730,1,L_SIZE),
				to_sfixed(0.9730,1,L_SIZE),
				to_sfixed(0.9730,1,L_SIZE),
				to_sfixed(0.9730,1,L_SIZE),
				to_sfixed(0.9730,1,L_SIZE),
				to_sfixed(0.9731,1,L_SIZE),
				to_sfixed(0.9731,1,L_SIZE),
				to_sfixed(0.9731,1,L_SIZE),
				to_sfixed(0.9731,1,L_SIZE),
				to_sfixed(0.9731,1,L_SIZE),
				to_sfixed(0.9731,1,L_SIZE),
				to_sfixed(0.9732,1,L_SIZE),
				to_sfixed(0.9732,1,L_SIZE),
				to_sfixed(0.9732,1,L_SIZE),
				to_sfixed(0.9732,1,L_SIZE),
				to_sfixed(0.9732,1,L_SIZE),
				to_sfixed(0.9733,1,L_SIZE),
				to_sfixed(0.9733,1,L_SIZE),
				to_sfixed(0.9733,1,L_SIZE),
				to_sfixed(0.9733,1,L_SIZE),
				to_sfixed(0.9733,1,L_SIZE),
				to_sfixed(0.9734,1,L_SIZE),
				to_sfixed(0.9734,1,L_SIZE),
				to_sfixed(0.9734,1,L_SIZE),
				to_sfixed(0.9734,1,L_SIZE),
				to_sfixed(0.9734,1,L_SIZE),
				to_sfixed(0.9735,1,L_SIZE),
				to_sfixed(0.9735,1,L_SIZE),
				to_sfixed(0.9735,1,L_SIZE),
				to_sfixed(0.9735,1,L_SIZE),
				to_sfixed(0.9735,1,L_SIZE),
				to_sfixed(0.9736,1,L_SIZE),
				to_sfixed(0.9736,1,L_SIZE),
				to_sfixed(0.9736,1,L_SIZE),
				to_sfixed(0.9736,1,L_SIZE),
				to_sfixed(0.9736,1,L_SIZE),
				to_sfixed(0.9736,1,L_SIZE),
				to_sfixed(0.9737,1,L_SIZE),
				to_sfixed(0.9737,1,L_SIZE),
				to_sfixed(0.9737,1,L_SIZE),
				to_sfixed(0.9737,1,L_SIZE),
				to_sfixed(0.9737,1,L_SIZE),
				to_sfixed(0.9738,1,L_SIZE),
				to_sfixed(0.9738,1,L_SIZE),
				to_sfixed(0.9738,1,L_SIZE),
				to_sfixed(0.9738,1,L_SIZE),
				to_sfixed(0.9738,1,L_SIZE),
				to_sfixed(0.9739,1,L_SIZE),
				to_sfixed(0.9739,1,L_SIZE),
				to_sfixed(0.9739,1,L_SIZE),
				to_sfixed(0.9739,1,L_SIZE),
				to_sfixed(0.9739,1,L_SIZE),
				to_sfixed(0.9740,1,L_SIZE),
				to_sfixed(0.9740,1,L_SIZE),
				to_sfixed(0.9740,1,L_SIZE),
				to_sfixed(0.9740,1,L_SIZE),
				to_sfixed(0.9740,1,L_SIZE),
				to_sfixed(0.9740,1,L_SIZE),
				to_sfixed(0.9741,1,L_SIZE),
				to_sfixed(0.9741,1,L_SIZE),
				to_sfixed(0.9741,1,L_SIZE),
				to_sfixed(0.9741,1,L_SIZE),
				to_sfixed(0.9741,1,L_SIZE),
				to_sfixed(0.9742,1,L_SIZE),
				to_sfixed(0.9742,1,L_SIZE),
				to_sfixed(0.9742,1,L_SIZE),
				to_sfixed(0.9742,1,L_SIZE),
				to_sfixed(0.9742,1,L_SIZE),
				to_sfixed(0.9743,1,L_SIZE),
				to_sfixed(0.9743,1,L_SIZE),
				to_sfixed(0.9743,1,L_SIZE),
				to_sfixed(0.9743,1,L_SIZE),
				to_sfixed(0.9743,1,L_SIZE),
				to_sfixed(0.9743,1,L_SIZE),
				to_sfixed(0.9744,1,L_SIZE),
				to_sfixed(0.9744,1,L_SIZE),
				to_sfixed(0.9744,1,L_SIZE),
				to_sfixed(0.9744,1,L_SIZE),
				to_sfixed(0.9744,1,L_SIZE),
				to_sfixed(0.9745,1,L_SIZE),
				to_sfixed(0.9745,1,L_SIZE),
				to_sfixed(0.9745,1,L_SIZE),
				to_sfixed(0.9745,1,L_SIZE),
				to_sfixed(0.9745,1,L_SIZE),
				to_sfixed(0.9745,1,L_SIZE),
				to_sfixed(0.9746,1,L_SIZE),
				to_sfixed(0.9746,1,L_SIZE),
				to_sfixed(0.9746,1,L_SIZE),
				to_sfixed(0.9746,1,L_SIZE),
				to_sfixed(0.9746,1,L_SIZE),
				to_sfixed(0.9747,1,L_SIZE),
				to_sfixed(0.9747,1,L_SIZE),
				to_sfixed(0.9747,1,L_SIZE),
				to_sfixed(0.9747,1,L_SIZE),
				to_sfixed(0.9747,1,L_SIZE),
				to_sfixed(0.9748,1,L_SIZE),
				to_sfixed(0.9748,1,L_SIZE),
				to_sfixed(0.9748,1,L_SIZE),
				to_sfixed(0.9748,1,L_SIZE),
				to_sfixed(0.9748,1,L_SIZE),
				to_sfixed(0.9748,1,L_SIZE),
				to_sfixed(0.9749,1,L_SIZE),
				to_sfixed(0.9749,1,L_SIZE),
				to_sfixed(0.9749,1,L_SIZE),
				to_sfixed(0.9749,1,L_SIZE),
				to_sfixed(0.9749,1,L_SIZE),
				to_sfixed(0.9750,1,L_SIZE),
				to_sfixed(0.9750,1,L_SIZE),
				to_sfixed(0.9750,1,L_SIZE),
				to_sfixed(0.9750,1,L_SIZE),
				to_sfixed(0.9750,1,L_SIZE),
				to_sfixed(0.9750,1,L_SIZE),
				to_sfixed(0.9751,1,L_SIZE),
				to_sfixed(0.9751,1,L_SIZE),
				to_sfixed(0.9751,1,L_SIZE),
				to_sfixed(0.9751,1,L_SIZE),
				to_sfixed(0.9751,1,L_SIZE),
				to_sfixed(0.9751,1,L_SIZE),
				to_sfixed(0.9752,1,L_SIZE),
				to_sfixed(0.9752,1,L_SIZE),
				to_sfixed(0.9752,1,L_SIZE),
				to_sfixed(0.9752,1,L_SIZE),
				to_sfixed(0.9752,1,L_SIZE),
				to_sfixed(0.9753,1,L_SIZE),
				to_sfixed(0.9753,1,L_SIZE),
				to_sfixed(0.9753,1,L_SIZE),
				to_sfixed(0.9753,1,L_SIZE),
				to_sfixed(0.9753,1,L_SIZE),
				to_sfixed(0.9753,1,L_SIZE),
				to_sfixed(0.9754,1,L_SIZE),
				to_sfixed(0.9754,1,L_SIZE),
				to_sfixed(0.9754,1,L_SIZE),
				to_sfixed(0.9754,1,L_SIZE),
				to_sfixed(0.9754,1,L_SIZE),
				to_sfixed(0.9755,1,L_SIZE),
				to_sfixed(0.9755,1,L_SIZE),
				to_sfixed(0.9755,1,L_SIZE),
				to_sfixed(0.9755,1,L_SIZE),
				to_sfixed(0.9755,1,L_SIZE),
				to_sfixed(0.9755,1,L_SIZE),
				to_sfixed(0.9756,1,L_SIZE),
				to_sfixed(0.9756,1,L_SIZE),
				to_sfixed(0.9756,1,L_SIZE),
				to_sfixed(0.9756,1,L_SIZE),
				to_sfixed(0.9756,1,L_SIZE),
				to_sfixed(0.9756,1,L_SIZE),
				to_sfixed(0.9757,1,L_SIZE),
				to_sfixed(0.9757,1,L_SIZE),
				to_sfixed(0.9757,1,L_SIZE),
				to_sfixed(0.9757,1,L_SIZE),
				to_sfixed(0.9757,1,L_SIZE),
				to_sfixed(0.9758,1,L_SIZE),
				to_sfixed(0.9758,1,L_SIZE),
				to_sfixed(0.9758,1,L_SIZE),
				to_sfixed(0.9758,1,L_SIZE),
				to_sfixed(0.9758,1,L_SIZE),
				to_sfixed(0.9758,1,L_SIZE),
				to_sfixed(0.9759,1,L_SIZE),
				to_sfixed(0.9759,1,L_SIZE),
				to_sfixed(0.9759,1,L_SIZE),
				to_sfixed(0.9759,1,L_SIZE),
				to_sfixed(0.9759,1,L_SIZE),
				to_sfixed(0.9759,1,L_SIZE),
				to_sfixed(0.9760,1,L_SIZE),
				to_sfixed(0.9760,1,L_SIZE),
				to_sfixed(0.9760,1,L_SIZE),
				to_sfixed(0.9760,1,L_SIZE),
				to_sfixed(0.9760,1,L_SIZE),
				to_sfixed(0.9760,1,L_SIZE),
				to_sfixed(0.9761,1,L_SIZE),
				to_sfixed(0.9761,1,L_SIZE),
				to_sfixed(0.9761,1,L_SIZE),
				to_sfixed(0.9761,1,L_SIZE),
				to_sfixed(0.9761,1,L_SIZE),
				to_sfixed(0.9762,1,L_SIZE),
				to_sfixed(0.9762,1,L_SIZE),
				to_sfixed(0.9762,1,L_SIZE),
				to_sfixed(0.9762,1,L_SIZE),
				to_sfixed(0.9762,1,L_SIZE),
				to_sfixed(0.9762,1,L_SIZE),
				to_sfixed(0.9763,1,L_SIZE),
				to_sfixed(0.9763,1,L_SIZE),
				to_sfixed(0.9763,1,L_SIZE),
				to_sfixed(0.9763,1,L_SIZE),
				to_sfixed(0.9763,1,L_SIZE),
				to_sfixed(0.9763,1,L_SIZE),
				to_sfixed(0.9764,1,L_SIZE),
				to_sfixed(0.9764,1,L_SIZE),
				to_sfixed(0.9764,1,L_SIZE),
				to_sfixed(0.9764,1,L_SIZE),
				to_sfixed(0.9764,1,L_SIZE),
				to_sfixed(0.9764,1,L_SIZE),
				to_sfixed(0.9765,1,L_SIZE),
				to_sfixed(0.9765,1,L_SIZE),
				to_sfixed(0.9765,1,L_SIZE),
				to_sfixed(0.9765,1,L_SIZE),
				to_sfixed(0.9765,1,L_SIZE),
				to_sfixed(0.9765,1,L_SIZE),
				to_sfixed(0.9766,1,L_SIZE),
				to_sfixed(0.9766,1,L_SIZE),
				to_sfixed(0.9766,1,L_SIZE),
				to_sfixed(0.9766,1,L_SIZE),
				to_sfixed(0.9766,1,L_SIZE),
				to_sfixed(0.9766,1,L_SIZE),
				to_sfixed(0.9767,1,L_SIZE),
				to_sfixed(0.9767,1,L_SIZE),
				to_sfixed(0.9767,1,L_SIZE),
				to_sfixed(0.9767,1,L_SIZE),
				to_sfixed(0.9767,1,L_SIZE),
				to_sfixed(0.9767,1,L_SIZE),
				to_sfixed(0.9768,1,L_SIZE),
				to_sfixed(0.9768,1,L_SIZE),
				to_sfixed(0.9768,1,L_SIZE),
				to_sfixed(0.9768,1,L_SIZE),
				to_sfixed(0.9768,1,L_SIZE),
				to_sfixed(0.9769,1,L_SIZE),
				to_sfixed(0.9769,1,L_SIZE),
				to_sfixed(0.9769,1,L_SIZE),
				to_sfixed(0.9769,1,L_SIZE),
				to_sfixed(0.9769,1,L_SIZE),
				to_sfixed(0.9769,1,L_SIZE),
				to_sfixed(0.9770,1,L_SIZE),
				to_sfixed(0.9770,1,L_SIZE),
				to_sfixed(0.9770,1,L_SIZE),
				to_sfixed(0.9770,1,L_SIZE),
				to_sfixed(0.9770,1,L_SIZE),
				to_sfixed(0.9770,1,L_SIZE),
				to_sfixed(0.9771,1,L_SIZE),
				to_sfixed(0.9771,1,L_SIZE),
				to_sfixed(0.9771,1,L_SIZE),
				to_sfixed(0.9771,1,L_SIZE),
				to_sfixed(0.9771,1,L_SIZE),
				to_sfixed(0.9771,1,L_SIZE),
				to_sfixed(0.9771,1,L_SIZE),
				to_sfixed(0.9772,1,L_SIZE),
				to_sfixed(0.9772,1,L_SIZE),
				to_sfixed(0.9772,1,L_SIZE),
				to_sfixed(0.9772,1,L_SIZE),
				to_sfixed(0.9772,1,L_SIZE),
				to_sfixed(0.9772,1,L_SIZE),
				to_sfixed(0.9773,1,L_SIZE),
				to_sfixed(0.9773,1,L_SIZE),
				to_sfixed(0.9773,1,L_SIZE),
				to_sfixed(0.9773,1,L_SIZE),
				to_sfixed(0.9773,1,L_SIZE),
				to_sfixed(0.9773,1,L_SIZE),
				to_sfixed(0.9774,1,L_SIZE),
				to_sfixed(0.9774,1,L_SIZE),
				to_sfixed(0.9774,1,L_SIZE),
				to_sfixed(0.9774,1,L_SIZE),
				to_sfixed(0.9774,1,L_SIZE),
				to_sfixed(0.9774,1,L_SIZE),
				to_sfixed(0.9775,1,L_SIZE),
				to_sfixed(0.9775,1,L_SIZE),
				to_sfixed(0.9775,1,L_SIZE),
				to_sfixed(0.9775,1,L_SIZE),
				to_sfixed(0.9775,1,L_SIZE),
				to_sfixed(0.9775,1,L_SIZE),
				to_sfixed(0.9776,1,L_SIZE),
				to_sfixed(0.9776,1,L_SIZE),
				to_sfixed(0.9776,1,L_SIZE),
				to_sfixed(0.9776,1,L_SIZE),
				to_sfixed(0.9776,1,L_SIZE),
				to_sfixed(0.9776,1,L_SIZE),
				to_sfixed(0.9777,1,L_SIZE),
				to_sfixed(0.9777,1,L_SIZE),
				to_sfixed(0.9777,1,L_SIZE),
				to_sfixed(0.9777,1,L_SIZE),
				to_sfixed(0.9777,1,L_SIZE),
				to_sfixed(0.9777,1,L_SIZE),
				to_sfixed(0.9778,1,L_SIZE),
				to_sfixed(0.9778,1,L_SIZE),
				to_sfixed(0.9778,1,L_SIZE),
				to_sfixed(0.9778,1,L_SIZE),
				to_sfixed(0.9778,1,L_SIZE),
				to_sfixed(0.9778,1,L_SIZE),
				to_sfixed(0.9779,1,L_SIZE),
				to_sfixed(0.9779,1,L_SIZE),
				to_sfixed(0.9779,1,L_SIZE),
				to_sfixed(0.9779,1,L_SIZE),
				to_sfixed(0.9779,1,L_SIZE),
				to_sfixed(0.9779,1,L_SIZE),
				to_sfixed(0.9779,1,L_SIZE),
				to_sfixed(0.9780,1,L_SIZE),
				to_sfixed(0.9780,1,L_SIZE),
				to_sfixed(0.9780,1,L_SIZE),
				to_sfixed(0.9780,1,L_SIZE),
				to_sfixed(0.9780,1,L_SIZE),
				to_sfixed(0.9780,1,L_SIZE),
				to_sfixed(0.9781,1,L_SIZE),
				to_sfixed(0.9781,1,L_SIZE),
				to_sfixed(0.9781,1,L_SIZE),
				to_sfixed(0.9781,1,L_SIZE),
				to_sfixed(0.9781,1,L_SIZE),
				to_sfixed(0.9781,1,L_SIZE),
				to_sfixed(0.9782,1,L_SIZE),
				to_sfixed(0.9782,1,L_SIZE),
				to_sfixed(0.9782,1,L_SIZE),
				to_sfixed(0.9782,1,L_SIZE),
				to_sfixed(0.9782,1,L_SIZE),
				to_sfixed(0.9782,1,L_SIZE),
				to_sfixed(0.9782,1,L_SIZE),
				to_sfixed(0.9783,1,L_SIZE),
				to_sfixed(0.9783,1,L_SIZE),
				to_sfixed(0.9783,1,L_SIZE),
				to_sfixed(0.9783,1,L_SIZE),
				to_sfixed(0.9783,1,L_SIZE),
				to_sfixed(0.9783,1,L_SIZE),
				to_sfixed(0.9784,1,L_SIZE),
				to_sfixed(0.9784,1,L_SIZE),
				to_sfixed(0.9784,1,L_SIZE),
				to_sfixed(0.9784,1,L_SIZE),
				to_sfixed(0.9784,1,L_SIZE),
				to_sfixed(0.9784,1,L_SIZE),
				to_sfixed(0.9785,1,L_SIZE),
				to_sfixed(0.9785,1,L_SIZE),
				to_sfixed(0.9785,1,L_SIZE),
				to_sfixed(0.9785,1,L_SIZE),
				to_sfixed(0.9785,1,L_SIZE),
				to_sfixed(0.9785,1,L_SIZE),
				to_sfixed(0.9785,1,L_SIZE),
				to_sfixed(0.9786,1,L_SIZE),
				to_sfixed(0.9786,1,L_SIZE),
				to_sfixed(0.9786,1,L_SIZE),
				to_sfixed(0.9786,1,L_SIZE),
				to_sfixed(0.9786,1,L_SIZE),
				to_sfixed(0.9786,1,L_SIZE),
				to_sfixed(0.9787,1,L_SIZE),
				to_sfixed(0.9787,1,L_SIZE),
				to_sfixed(0.9787,1,L_SIZE),
				to_sfixed(0.9787,1,L_SIZE),
				to_sfixed(0.9787,1,L_SIZE),
				to_sfixed(0.9787,1,L_SIZE),
				to_sfixed(0.9787,1,L_SIZE),
				to_sfixed(0.9788,1,L_SIZE),
				to_sfixed(0.9788,1,L_SIZE),
				to_sfixed(0.9788,1,L_SIZE),
				to_sfixed(0.9788,1,L_SIZE),
				to_sfixed(0.9788,1,L_SIZE),
				to_sfixed(0.9788,1,L_SIZE),
				to_sfixed(0.9789,1,L_SIZE),
				to_sfixed(0.9789,1,L_SIZE),
				to_sfixed(0.9789,1,L_SIZE),
				to_sfixed(0.9789,1,L_SIZE),
				to_sfixed(0.9789,1,L_SIZE),
				to_sfixed(0.9789,1,L_SIZE),
				to_sfixed(0.9789,1,L_SIZE),
				to_sfixed(0.9790,1,L_SIZE),
				to_sfixed(0.9790,1,L_SIZE),
				to_sfixed(0.9790,1,L_SIZE),
				to_sfixed(0.9790,1,L_SIZE),
				to_sfixed(0.9790,1,L_SIZE),
				to_sfixed(0.9790,1,L_SIZE),
				to_sfixed(0.9791,1,L_SIZE),
				to_sfixed(0.9791,1,L_SIZE),
				to_sfixed(0.9791,1,L_SIZE),
				to_sfixed(0.9791,1,L_SIZE),
				to_sfixed(0.9791,1,L_SIZE),
				to_sfixed(0.9791,1,L_SIZE),
				to_sfixed(0.9791,1,L_SIZE),
				to_sfixed(0.9792,1,L_SIZE),
				to_sfixed(0.9792,1,L_SIZE),
				to_sfixed(0.9792,1,L_SIZE),
				to_sfixed(0.9792,1,L_SIZE),
				to_sfixed(0.9792,1,L_SIZE),
				to_sfixed(0.9792,1,L_SIZE),
				to_sfixed(0.9792,1,L_SIZE),
				to_sfixed(0.9793,1,L_SIZE),
				to_sfixed(0.9793,1,L_SIZE),
				to_sfixed(0.9793,1,L_SIZE),
				to_sfixed(0.9793,1,L_SIZE),
				to_sfixed(0.9793,1,L_SIZE),
				to_sfixed(0.9793,1,L_SIZE),
				to_sfixed(0.9794,1,L_SIZE),
				to_sfixed(0.9794,1,L_SIZE),
				to_sfixed(0.9794,1,L_SIZE),
				to_sfixed(0.9794,1,L_SIZE),
				to_sfixed(0.9794,1,L_SIZE),
				to_sfixed(0.9794,1,L_SIZE),
				to_sfixed(0.9794,1,L_SIZE),
				to_sfixed(0.9795,1,L_SIZE),
				to_sfixed(0.9795,1,L_SIZE),
				to_sfixed(0.9795,1,L_SIZE),
				to_sfixed(0.9795,1,L_SIZE),
				to_sfixed(0.9795,1,L_SIZE),
				to_sfixed(0.9795,1,L_SIZE),
				to_sfixed(0.9795,1,L_SIZE),
				to_sfixed(0.9796,1,L_SIZE),
				to_sfixed(0.9796,1,L_SIZE),
				to_sfixed(0.9796,1,L_SIZE),
				to_sfixed(0.9796,1,L_SIZE),
				to_sfixed(0.9796,1,L_SIZE),
				to_sfixed(0.9796,1,L_SIZE),
				to_sfixed(0.9797,1,L_SIZE),
				to_sfixed(0.9797,1,L_SIZE),
				to_sfixed(0.9797,1,L_SIZE),
				to_sfixed(0.9797,1,L_SIZE),
				to_sfixed(0.9797,1,L_SIZE),
				to_sfixed(0.9797,1,L_SIZE),
				to_sfixed(0.9797,1,L_SIZE),
				to_sfixed(0.9798,1,L_SIZE),
				to_sfixed(0.9798,1,L_SIZE),
				to_sfixed(0.9798,1,L_SIZE),
				to_sfixed(0.9798,1,L_SIZE),
				to_sfixed(0.9798,1,L_SIZE),
				to_sfixed(0.9798,1,L_SIZE),
				to_sfixed(0.9798,1,L_SIZE),
				to_sfixed(0.9799,1,L_SIZE),
				to_sfixed(0.9799,1,L_SIZE),
				to_sfixed(0.9799,1,L_SIZE),
				to_sfixed(0.9799,1,L_SIZE),
				to_sfixed(0.9799,1,L_SIZE),
				to_sfixed(0.9799,1,L_SIZE),
				to_sfixed(0.9799,1,L_SIZE),
				to_sfixed(0.9800,1,L_SIZE),
				to_sfixed(0.9800,1,L_SIZE),
				to_sfixed(0.9800,1,L_SIZE),
				to_sfixed(0.9800,1,L_SIZE),
				to_sfixed(0.9800,1,L_SIZE),
				to_sfixed(0.9800,1,L_SIZE),
				to_sfixed(0.9800,1,L_SIZE),
				to_sfixed(0.9801,1,L_SIZE),
				to_sfixed(0.9801,1,L_SIZE),
				to_sfixed(0.9801,1,L_SIZE),
				to_sfixed(0.9801,1,L_SIZE),
				to_sfixed(0.9801,1,L_SIZE),
				to_sfixed(0.9801,1,L_SIZE),
				to_sfixed(0.9801,1,L_SIZE),
				to_sfixed(0.9802,1,L_SIZE),
				to_sfixed(0.9802,1,L_SIZE),
				to_sfixed(0.9802,1,L_SIZE),
				to_sfixed(0.9802,1,L_SIZE),
				to_sfixed(0.9802,1,L_SIZE),
				to_sfixed(0.9802,1,L_SIZE),
				to_sfixed(0.9802,1,L_SIZE),
				to_sfixed(0.9803,1,L_SIZE),
				to_sfixed(0.9803,1,L_SIZE),
				to_sfixed(0.9803,1,L_SIZE),
				to_sfixed(0.9803,1,L_SIZE),
				to_sfixed(0.9803,1,L_SIZE),
				to_sfixed(0.9803,1,L_SIZE),
				to_sfixed(0.9803,1,L_SIZE),
				to_sfixed(0.9804,1,L_SIZE),
				to_sfixed(0.9804,1,L_SIZE),
				to_sfixed(0.9804,1,L_SIZE),
				to_sfixed(0.9804,1,L_SIZE),
				to_sfixed(0.9804,1,L_SIZE),
				to_sfixed(0.9804,1,L_SIZE),
				to_sfixed(0.9804,1,L_SIZE),
				to_sfixed(0.9805,1,L_SIZE),
				to_sfixed(0.9805,1,L_SIZE),
				to_sfixed(0.9805,1,L_SIZE),
				to_sfixed(0.9805,1,L_SIZE),
				to_sfixed(0.9805,1,L_SIZE),
				to_sfixed(0.9805,1,L_SIZE),
				to_sfixed(0.9805,1,L_SIZE),
				to_sfixed(0.9806,1,L_SIZE),
				to_sfixed(0.9806,1,L_SIZE),
				to_sfixed(0.9806,1,L_SIZE),
				to_sfixed(0.9806,1,L_SIZE),
				to_sfixed(0.9806,1,L_SIZE),
				to_sfixed(0.9806,1,L_SIZE),
				to_sfixed(0.9806,1,L_SIZE),
				to_sfixed(0.9807,1,L_SIZE),
				to_sfixed(0.9807,1,L_SIZE),
				to_sfixed(0.9807,1,L_SIZE),
				to_sfixed(0.9807,1,L_SIZE),
				to_sfixed(0.9807,1,L_SIZE),
				to_sfixed(0.9807,1,L_SIZE),
				to_sfixed(0.9807,1,L_SIZE),
				to_sfixed(0.9808,1,L_SIZE),
				to_sfixed(0.9808,1,L_SIZE),
				to_sfixed(0.9808,1,L_SIZE),
				to_sfixed(0.9808,1,L_SIZE),
				to_sfixed(0.9808,1,L_SIZE),
				to_sfixed(0.9808,1,L_SIZE),
				to_sfixed(0.9808,1,L_SIZE),
				to_sfixed(0.9809,1,L_SIZE),
				to_sfixed(0.9809,1,L_SIZE),
				to_sfixed(0.9809,1,L_SIZE),
				to_sfixed(0.9809,1,L_SIZE),
				to_sfixed(0.9809,1,L_SIZE),
				to_sfixed(0.9809,1,L_SIZE),
				to_sfixed(0.9809,1,L_SIZE),
				to_sfixed(0.9810,1,L_SIZE),
				to_sfixed(0.9810,1,L_SIZE),
				to_sfixed(0.9810,1,L_SIZE),
				to_sfixed(0.9810,1,L_SIZE),
				to_sfixed(0.9810,1,L_SIZE),
				to_sfixed(0.9810,1,L_SIZE),
				to_sfixed(0.9810,1,L_SIZE),
				to_sfixed(0.9810,1,L_SIZE),
				to_sfixed(0.9811,1,L_SIZE),
				to_sfixed(0.9811,1,L_SIZE),
				to_sfixed(0.9811,1,L_SIZE),
				to_sfixed(0.9811,1,L_SIZE),
				to_sfixed(0.9811,1,L_SIZE),
				to_sfixed(0.9811,1,L_SIZE),
				to_sfixed(0.9811,1,L_SIZE),
				to_sfixed(0.9812,1,L_SIZE),
				to_sfixed(0.9812,1,L_SIZE),
				to_sfixed(0.9812,1,L_SIZE),
				to_sfixed(0.9812,1,L_SIZE),
				to_sfixed(0.9812,1,L_SIZE),
				to_sfixed(0.9812,1,L_SIZE),
				to_sfixed(0.9812,1,L_SIZE),
				to_sfixed(0.9813,1,L_SIZE),
				to_sfixed(0.9813,1,L_SIZE),
				to_sfixed(0.9813,1,L_SIZE),
				to_sfixed(0.9813,1,L_SIZE),
				to_sfixed(0.9813,1,L_SIZE),
				to_sfixed(0.9813,1,L_SIZE),
				to_sfixed(0.9813,1,L_SIZE),
				to_sfixed(0.9813,1,L_SIZE),
				to_sfixed(0.9814,1,L_SIZE),
				to_sfixed(0.9814,1,L_SIZE),
				to_sfixed(0.9814,1,L_SIZE),
				to_sfixed(0.9814,1,L_SIZE),
				to_sfixed(0.9814,1,L_SIZE),
				to_sfixed(0.9814,1,L_SIZE),
				to_sfixed(0.9814,1,L_SIZE),
				to_sfixed(0.9815,1,L_SIZE),
				to_sfixed(0.9815,1,L_SIZE),
				to_sfixed(0.9815,1,L_SIZE),
				to_sfixed(0.9815,1,L_SIZE),
				to_sfixed(0.9815,1,L_SIZE),
				to_sfixed(0.9815,1,L_SIZE),
				to_sfixed(0.9815,1,L_SIZE),
				to_sfixed(0.9815,1,L_SIZE),
				to_sfixed(0.9816,1,L_SIZE),
				to_sfixed(0.9816,1,L_SIZE),
				to_sfixed(0.9816,1,L_SIZE),
				to_sfixed(0.9816,1,L_SIZE),
				to_sfixed(0.9816,1,L_SIZE),
				to_sfixed(0.9816,1,L_SIZE),
				to_sfixed(0.9816,1,L_SIZE),
				to_sfixed(0.9817,1,L_SIZE),
				to_sfixed(0.9817,1,L_SIZE),
				to_sfixed(0.9817,1,L_SIZE),
				to_sfixed(0.9817,1,L_SIZE),
				to_sfixed(0.9817,1,L_SIZE),
				to_sfixed(0.9817,1,L_SIZE),
				to_sfixed(0.9817,1,L_SIZE),
				to_sfixed(0.9817,1,L_SIZE),
				to_sfixed(0.9818,1,L_SIZE),
				to_sfixed(0.9818,1,L_SIZE),
				to_sfixed(0.9818,1,L_SIZE),
				to_sfixed(0.9818,1,L_SIZE),
				to_sfixed(0.9818,1,L_SIZE),
				to_sfixed(0.9818,1,L_SIZE),
				to_sfixed(0.9818,1,L_SIZE),
				to_sfixed(0.9819,1,L_SIZE),
				to_sfixed(0.9819,1,L_SIZE),
				to_sfixed(0.9819,1,L_SIZE),
				to_sfixed(0.9819,1,L_SIZE),
				to_sfixed(0.9819,1,L_SIZE),
				to_sfixed(0.9819,1,L_SIZE),
				to_sfixed(0.9819,1,L_SIZE),
				to_sfixed(0.9819,1,L_SIZE),
				to_sfixed(0.9820,1,L_SIZE),
				to_sfixed(0.9820,1,L_SIZE),
				to_sfixed(0.9820,1,L_SIZE),
				to_sfixed(0.9820,1,L_SIZE),
				to_sfixed(0.9820,1,L_SIZE),
				to_sfixed(0.9820,1,L_SIZE),
				to_sfixed(0.9820,1,L_SIZE),
				to_sfixed(0.9821,1,L_SIZE),
				to_sfixed(0.9821,1,L_SIZE),
				to_sfixed(0.9821,1,L_SIZE),
				to_sfixed(0.9821,1,L_SIZE),
				to_sfixed(0.9821,1,L_SIZE),
				to_sfixed(0.9821,1,L_SIZE),
				to_sfixed(0.9821,1,L_SIZE),
				to_sfixed(0.9821,1,L_SIZE),
				to_sfixed(0.9822,1,L_SIZE),
				to_sfixed(0.9822,1,L_SIZE),
				to_sfixed(0.9822,1,L_SIZE),
				to_sfixed(0.9822,1,L_SIZE),
				to_sfixed(0.9822,1,L_SIZE),
				to_sfixed(0.9822,1,L_SIZE),
				to_sfixed(0.9822,1,L_SIZE),
				to_sfixed(0.9822,1,L_SIZE),
				to_sfixed(0.9823,1,L_SIZE),
				to_sfixed(0.9823,1,L_SIZE),
				to_sfixed(0.9823,1,L_SIZE),
				to_sfixed(0.9823,1,L_SIZE),
				to_sfixed(0.9823,1,L_SIZE),
				to_sfixed(0.9823,1,L_SIZE),
				to_sfixed(0.9823,1,L_SIZE),
				to_sfixed(0.9823,1,L_SIZE),
				to_sfixed(0.9824,1,L_SIZE),
				to_sfixed(0.9824,1,L_SIZE),
				to_sfixed(0.9824,1,L_SIZE),
				to_sfixed(0.9824,1,L_SIZE),
				to_sfixed(0.9824,1,L_SIZE),
				to_sfixed(0.9824,1,L_SIZE),
				to_sfixed(0.9824,1,L_SIZE),
				to_sfixed(0.9825,1,L_SIZE),
				to_sfixed(0.9825,1,L_SIZE),
				to_sfixed(0.9825,1,L_SIZE),
				to_sfixed(0.9825,1,L_SIZE),
				to_sfixed(0.9825,1,L_SIZE),
				to_sfixed(0.9825,1,L_SIZE),
				to_sfixed(0.9825,1,L_SIZE),
				to_sfixed(0.9825,1,L_SIZE),
				to_sfixed(0.9826,1,L_SIZE),
				to_sfixed(0.9826,1,L_SIZE),
				to_sfixed(0.9826,1,L_SIZE),
				to_sfixed(0.9826,1,L_SIZE),
				to_sfixed(0.9826,1,L_SIZE),
				to_sfixed(0.9826,1,L_SIZE),
				to_sfixed(0.9826,1,L_SIZE),
				to_sfixed(0.9826,1,L_SIZE),
				to_sfixed(0.9827,1,L_SIZE),
				to_sfixed(0.9827,1,L_SIZE),
				to_sfixed(0.9827,1,L_SIZE),
				to_sfixed(0.9827,1,L_SIZE),
				to_sfixed(0.9827,1,L_SIZE),
				to_sfixed(0.9827,1,L_SIZE),
				to_sfixed(0.9827,1,L_SIZE),
				to_sfixed(0.9827,1,L_SIZE),
				to_sfixed(0.9828,1,L_SIZE),
				to_sfixed(0.9828,1,L_SIZE),
				to_sfixed(0.9828,1,L_SIZE),
				to_sfixed(0.9828,1,L_SIZE),
				to_sfixed(0.9828,1,L_SIZE),
				to_sfixed(0.9828,1,L_SIZE),
				to_sfixed(0.9828,1,L_SIZE),
				to_sfixed(0.9828,1,L_SIZE),
				to_sfixed(0.9829,1,L_SIZE),
				to_sfixed(0.9829,1,L_SIZE),
				to_sfixed(0.9829,1,L_SIZE),
				to_sfixed(0.9829,1,L_SIZE),
				to_sfixed(0.9829,1,L_SIZE),
				to_sfixed(0.9829,1,L_SIZE),
				to_sfixed(0.9829,1,L_SIZE),
				to_sfixed(0.9829,1,L_SIZE),
				to_sfixed(0.9830,1,L_SIZE),
				to_sfixed(0.9830,1,L_SIZE),
				to_sfixed(0.9830,1,L_SIZE),
				to_sfixed(0.9830,1,L_SIZE),
				to_sfixed(0.9830,1,L_SIZE),
				to_sfixed(0.9830,1,L_SIZE),
				to_sfixed(0.9830,1,L_SIZE),
				to_sfixed(0.9830,1,L_SIZE),
				to_sfixed(0.9831,1,L_SIZE),
				to_sfixed(0.9831,1,L_SIZE),
				to_sfixed(0.9831,1,L_SIZE),
				to_sfixed(0.9831,1,L_SIZE),
				to_sfixed(0.9831,1,L_SIZE),
				to_sfixed(0.9831,1,L_SIZE),
				to_sfixed(0.9831,1,L_SIZE),
				to_sfixed(0.9831,1,L_SIZE),
				to_sfixed(0.9831,1,L_SIZE),
				to_sfixed(0.9832,1,L_SIZE),
				to_sfixed(0.9832,1,L_SIZE),
				to_sfixed(0.9832,1,L_SIZE),
				to_sfixed(0.9832,1,L_SIZE),
				to_sfixed(0.9832,1,L_SIZE),
				to_sfixed(0.9832,1,L_SIZE),
				to_sfixed(0.9832,1,L_SIZE),
				to_sfixed(0.9832,1,L_SIZE),
				to_sfixed(0.9833,1,L_SIZE),
				to_sfixed(0.9833,1,L_SIZE),
				to_sfixed(0.9833,1,L_SIZE),
				to_sfixed(0.9833,1,L_SIZE),
				to_sfixed(0.9833,1,L_SIZE),
				to_sfixed(0.9833,1,L_SIZE),
				to_sfixed(0.9833,1,L_SIZE),
				to_sfixed(0.9833,1,L_SIZE),
				to_sfixed(0.9834,1,L_SIZE),
				to_sfixed(0.9834,1,L_SIZE),
				to_sfixed(0.9834,1,L_SIZE),
				to_sfixed(0.9834,1,L_SIZE),
				to_sfixed(0.9834,1,L_SIZE),
				to_sfixed(0.9834,1,L_SIZE),
				to_sfixed(0.9834,1,L_SIZE),
				to_sfixed(0.9834,1,L_SIZE),
				to_sfixed(0.9835,1,L_SIZE),
				to_sfixed(0.9835,1,L_SIZE),
				to_sfixed(0.9835,1,L_SIZE),
				to_sfixed(0.9835,1,L_SIZE),
				to_sfixed(0.9835,1,L_SIZE),
				to_sfixed(0.9835,1,L_SIZE),
				to_sfixed(0.9835,1,L_SIZE),
				to_sfixed(0.9835,1,L_SIZE),
				to_sfixed(0.9835,1,L_SIZE),
				to_sfixed(0.9836,1,L_SIZE),
				to_sfixed(0.9836,1,L_SIZE),
				to_sfixed(0.9836,1,L_SIZE),
				to_sfixed(0.9836,1,L_SIZE),
				to_sfixed(0.9836,1,L_SIZE),
				to_sfixed(0.9836,1,L_SIZE),
				to_sfixed(0.9836,1,L_SIZE),
				to_sfixed(0.9836,1,L_SIZE),
				to_sfixed(0.9837,1,L_SIZE),
				to_sfixed(0.9837,1,L_SIZE),
				to_sfixed(0.9837,1,L_SIZE),
				to_sfixed(0.9837,1,L_SIZE),
				to_sfixed(0.9837,1,L_SIZE),
				to_sfixed(0.9837,1,L_SIZE),
				to_sfixed(0.9837,1,L_SIZE),
				to_sfixed(0.9837,1,L_SIZE),
				to_sfixed(0.9838,1,L_SIZE),
				to_sfixed(0.9838,1,L_SIZE),
				to_sfixed(0.9838,1,L_SIZE),
				to_sfixed(0.9838,1,L_SIZE),
				to_sfixed(0.9838,1,L_SIZE),
				to_sfixed(0.9838,1,L_SIZE),
				to_sfixed(0.9838,1,L_SIZE),
				to_sfixed(0.9838,1,L_SIZE),
				to_sfixed(0.9838,1,L_SIZE),
				to_sfixed(0.9839,1,L_SIZE),
				to_sfixed(0.9839,1,L_SIZE),
				to_sfixed(0.9839,1,L_SIZE),
				to_sfixed(0.9839,1,L_SIZE),
				to_sfixed(0.9839,1,L_SIZE),
				to_sfixed(0.9839,1,L_SIZE),
				to_sfixed(0.9839,1,L_SIZE),
				to_sfixed(0.9839,1,L_SIZE),
				to_sfixed(0.9840,1,L_SIZE),
				to_sfixed(0.9840,1,L_SIZE),
				to_sfixed(0.9840,1,L_SIZE),
				to_sfixed(0.9840,1,L_SIZE),
				to_sfixed(0.9840,1,L_SIZE),
				to_sfixed(0.9840,1,L_SIZE),
				to_sfixed(0.9840,1,L_SIZE),
				to_sfixed(0.9840,1,L_SIZE),
				to_sfixed(0.9840,1,L_SIZE),
				to_sfixed(0.9841,1,L_SIZE),
				to_sfixed(0.9841,1,L_SIZE),
				to_sfixed(0.9841,1,L_SIZE),
				to_sfixed(0.9841,1,L_SIZE),
				to_sfixed(0.9841,1,L_SIZE),
				to_sfixed(0.9841,1,L_SIZE),
				to_sfixed(0.9841,1,L_SIZE),
				to_sfixed(0.9841,1,L_SIZE),
				to_sfixed(0.9841,1,L_SIZE),
				to_sfixed(0.9842,1,L_SIZE),
				to_sfixed(0.9842,1,L_SIZE),
				to_sfixed(0.9842,1,L_SIZE),
				to_sfixed(0.9842,1,L_SIZE),
				to_sfixed(0.9842,1,L_SIZE),
				to_sfixed(0.9842,1,L_SIZE),
				to_sfixed(0.9842,1,L_SIZE),
				to_sfixed(0.9842,1,L_SIZE),
				to_sfixed(0.9843,1,L_SIZE),
				to_sfixed(0.9843,1,L_SIZE),
				to_sfixed(0.9843,1,L_SIZE),
				to_sfixed(0.9843,1,L_SIZE),
				to_sfixed(0.9843,1,L_SIZE),
				to_sfixed(0.9843,1,L_SIZE),
				to_sfixed(0.9843,1,L_SIZE),
				to_sfixed(0.9843,1,L_SIZE),
				to_sfixed(0.9843,1,L_SIZE),
				to_sfixed(0.9844,1,L_SIZE),
				to_sfixed(0.9844,1,L_SIZE),
				to_sfixed(0.9844,1,L_SIZE),
				to_sfixed(0.9844,1,L_SIZE),
				to_sfixed(0.9844,1,L_SIZE),
				to_sfixed(0.9844,1,L_SIZE),
				to_sfixed(0.9844,1,L_SIZE),
				to_sfixed(0.9844,1,L_SIZE),
				to_sfixed(0.9844,1,L_SIZE),
				to_sfixed(0.9845,1,L_SIZE),
				to_sfixed(0.9845,1,L_SIZE),
				to_sfixed(0.9845,1,L_SIZE),
				to_sfixed(0.9845,1,L_SIZE),
				to_sfixed(0.9845,1,L_SIZE),
				to_sfixed(0.9845,1,L_SIZE),
				to_sfixed(0.9845,1,L_SIZE),
				to_sfixed(0.9845,1,L_SIZE),
				to_sfixed(0.9845,1,L_SIZE),
				to_sfixed(0.9846,1,L_SIZE),
				to_sfixed(0.9846,1,L_SIZE),
				to_sfixed(0.9846,1,L_SIZE),
				to_sfixed(0.9846,1,L_SIZE),
				to_sfixed(0.9846,1,L_SIZE),
				to_sfixed(0.9846,1,L_SIZE),
				to_sfixed(0.9846,1,L_SIZE),
				to_sfixed(0.9846,1,L_SIZE),
				to_sfixed(0.9846,1,L_SIZE),
				to_sfixed(0.9847,1,L_SIZE),
				to_sfixed(0.9847,1,L_SIZE),
				to_sfixed(0.9847,1,L_SIZE),
				to_sfixed(0.9847,1,L_SIZE),
				to_sfixed(0.9847,1,L_SIZE),
				to_sfixed(0.9847,1,L_SIZE),
				to_sfixed(0.9847,1,L_SIZE),
				to_sfixed(0.9847,1,L_SIZE),
				to_sfixed(0.9847,1,L_SIZE),
				to_sfixed(0.9848,1,L_SIZE),
				to_sfixed(0.9848,1,L_SIZE),
				to_sfixed(0.9848,1,L_SIZE),
				to_sfixed(0.9848,1,L_SIZE),
				to_sfixed(0.9848,1,L_SIZE),
				to_sfixed(0.9848,1,L_SIZE),
				to_sfixed(0.9848,1,L_SIZE),
				to_sfixed(0.9848,1,L_SIZE),
				to_sfixed(0.9848,1,L_SIZE),
				to_sfixed(0.9849,1,L_SIZE),
				to_sfixed(0.9849,1,L_SIZE),
				to_sfixed(0.9849,1,L_SIZE),
				to_sfixed(0.9849,1,L_SIZE),
				to_sfixed(0.9849,1,L_SIZE),
				to_sfixed(0.9849,1,L_SIZE),
				to_sfixed(0.9849,1,L_SIZE),
				to_sfixed(0.9849,1,L_SIZE),
				to_sfixed(0.9849,1,L_SIZE),
				to_sfixed(0.9850,1,L_SIZE),
				to_sfixed(0.9850,1,L_SIZE),
				to_sfixed(0.9850,1,L_SIZE),
				to_sfixed(0.9850,1,L_SIZE),
				to_sfixed(0.9850,1,L_SIZE),
				to_sfixed(0.9850,1,L_SIZE),
				to_sfixed(0.9850,1,L_SIZE),
				to_sfixed(0.9850,1,L_SIZE),
				to_sfixed(0.9850,1,L_SIZE),
				to_sfixed(0.9851,1,L_SIZE),
				to_sfixed(0.9851,1,L_SIZE),
				to_sfixed(0.9851,1,L_SIZE),
				to_sfixed(0.9851,1,L_SIZE),
				to_sfixed(0.9851,1,L_SIZE),
				to_sfixed(0.9851,1,L_SIZE),
				to_sfixed(0.9851,1,L_SIZE),
				to_sfixed(0.9851,1,L_SIZE),
				to_sfixed(0.9851,1,L_SIZE),
				to_sfixed(0.9852,1,L_SIZE),
				to_sfixed(0.9852,1,L_SIZE),
				to_sfixed(0.9852,1,L_SIZE),
				to_sfixed(0.9852,1,L_SIZE),
				to_sfixed(0.9852,1,L_SIZE),
				to_sfixed(0.9852,1,L_SIZE),
				to_sfixed(0.9852,1,L_SIZE),
				to_sfixed(0.9852,1,L_SIZE),
				to_sfixed(0.9852,1,L_SIZE),
				to_sfixed(0.9852,1,L_SIZE),
				to_sfixed(0.9853,1,L_SIZE),
				to_sfixed(0.9853,1,L_SIZE),
				to_sfixed(0.9853,1,L_SIZE),
				to_sfixed(0.9853,1,L_SIZE),
				to_sfixed(0.9853,1,L_SIZE),
				to_sfixed(0.9853,1,L_SIZE),
				to_sfixed(0.9853,1,L_SIZE),
				to_sfixed(0.9853,1,L_SIZE),
				to_sfixed(0.9853,1,L_SIZE),
				to_sfixed(0.9854,1,L_SIZE),
				to_sfixed(0.9854,1,L_SIZE),
				to_sfixed(0.9854,1,L_SIZE),
				to_sfixed(0.9854,1,L_SIZE),
				to_sfixed(0.9854,1,L_SIZE),
				to_sfixed(0.9854,1,L_SIZE),
				to_sfixed(0.9854,1,L_SIZE),
				to_sfixed(0.9854,1,L_SIZE),
				to_sfixed(0.9854,1,L_SIZE),
				to_sfixed(0.9855,1,L_SIZE),
				to_sfixed(0.9855,1,L_SIZE),
				to_sfixed(0.9855,1,L_SIZE),
				to_sfixed(0.9855,1,L_SIZE),
				to_sfixed(0.9855,1,L_SIZE),
				to_sfixed(0.9855,1,L_SIZE),
				to_sfixed(0.9855,1,L_SIZE),
				to_sfixed(0.9855,1,L_SIZE),
				to_sfixed(0.9855,1,L_SIZE),
				to_sfixed(0.9855,1,L_SIZE),
				to_sfixed(0.9856,1,L_SIZE),
				to_sfixed(0.9856,1,L_SIZE),
				to_sfixed(0.9856,1,L_SIZE),
				to_sfixed(0.9856,1,L_SIZE),
				to_sfixed(0.9856,1,L_SIZE),
				to_sfixed(0.9856,1,L_SIZE),
				to_sfixed(0.9856,1,L_SIZE),
				to_sfixed(0.9856,1,L_SIZE),
				to_sfixed(0.9856,1,L_SIZE),
				to_sfixed(0.9856,1,L_SIZE),
				to_sfixed(0.9857,1,L_SIZE),
				to_sfixed(0.9857,1,L_SIZE),
				to_sfixed(0.9857,1,L_SIZE),
				to_sfixed(0.9857,1,L_SIZE),
				to_sfixed(0.9857,1,L_SIZE),
				to_sfixed(0.9857,1,L_SIZE),
				to_sfixed(0.9857,1,L_SIZE),
				to_sfixed(0.9857,1,L_SIZE),
				to_sfixed(0.9857,1,L_SIZE),
				to_sfixed(0.9858,1,L_SIZE),
				to_sfixed(0.9858,1,L_SIZE),
				to_sfixed(0.9858,1,L_SIZE),
				to_sfixed(0.9858,1,L_SIZE),
				to_sfixed(0.9858,1,L_SIZE),
				to_sfixed(0.9858,1,L_SIZE),
				to_sfixed(0.9858,1,L_SIZE),
				to_sfixed(0.9858,1,L_SIZE),
				to_sfixed(0.9858,1,L_SIZE),
				to_sfixed(0.9858,1,L_SIZE),
				to_sfixed(0.9859,1,L_SIZE),
				to_sfixed(0.9859,1,L_SIZE),
				to_sfixed(0.9859,1,L_SIZE),
				to_sfixed(0.9859,1,L_SIZE),
				to_sfixed(0.9859,1,L_SIZE),
				to_sfixed(0.9859,1,L_SIZE),
				to_sfixed(0.9859,1,L_SIZE),
				to_sfixed(0.9859,1,L_SIZE),
				to_sfixed(0.9859,1,L_SIZE),
				to_sfixed(0.9859,1,L_SIZE),
				to_sfixed(0.9860,1,L_SIZE),
				to_sfixed(0.9860,1,L_SIZE),
				to_sfixed(0.9860,1,L_SIZE),
				to_sfixed(0.9860,1,L_SIZE),
				to_sfixed(0.9860,1,L_SIZE),
				to_sfixed(0.9860,1,L_SIZE),
				to_sfixed(0.9860,1,L_SIZE),
				to_sfixed(0.9860,1,L_SIZE),
				to_sfixed(0.9860,1,L_SIZE),
				to_sfixed(0.9861,1,L_SIZE),
				to_sfixed(0.9861,1,L_SIZE),
				to_sfixed(0.9861,1,L_SIZE),
				to_sfixed(0.9861,1,L_SIZE),
				to_sfixed(0.9861,1,L_SIZE),
				to_sfixed(0.9861,1,L_SIZE),
				to_sfixed(0.9861,1,L_SIZE),
				to_sfixed(0.9861,1,L_SIZE),
				to_sfixed(0.9861,1,L_SIZE),
				to_sfixed(0.9861,1,L_SIZE),
				to_sfixed(0.9862,1,L_SIZE),
				to_sfixed(0.9862,1,L_SIZE),
				to_sfixed(0.9862,1,L_SIZE),
				to_sfixed(0.9862,1,L_SIZE),
				to_sfixed(0.9862,1,L_SIZE),
				to_sfixed(0.9862,1,L_SIZE),
				to_sfixed(0.9862,1,L_SIZE),
				to_sfixed(0.9862,1,L_SIZE),
				to_sfixed(0.9862,1,L_SIZE),
				to_sfixed(0.9862,1,L_SIZE),
				to_sfixed(0.9863,1,L_SIZE),
				to_sfixed(0.9863,1,L_SIZE),
				to_sfixed(0.9863,1,L_SIZE),
				to_sfixed(0.9863,1,L_SIZE),
				to_sfixed(0.9863,1,L_SIZE),
				to_sfixed(0.9863,1,L_SIZE),
				to_sfixed(0.9863,1,L_SIZE),
				to_sfixed(0.9863,1,L_SIZE),
				to_sfixed(0.9863,1,L_SIZE),
				to_sfixed(0.9863,1,L_SIZE),
				to_sfixed(0.9864,1,L_SIZE),
				to_sfixed(0.9864,1,L_SIZE),
				to_sfixed(0.9864,1,L_SIZE),
				to_sfixed(0.9864,1,L_SIZE),
				to_sfixed(0.9864,1,L_SIZE),
				to_sfixed(0.9864,1,L_SIZE),
				to_sfixed(0.9864,1,L_SIZE),
				to_sfixed(0.9864,1,L_SIZE),
				to_sfixed(0.9864,1,L_SIZE),
				to_sfixed(0.9864,1,L_SIZE),
				to_sfixed(0.9865,1,L_SIZE),
				to_sfixed(0.9865,1,L_SIZE),
				to_sfixed(0.9865,1,L_SIZE),
				to_sfixed(0.9865,1,L_SIZE),
				to_sfixed(0.9865,1,L_SIZE),
				to_sfixed(0.9865,1,L_SIZE),
				to_sfixed(0.9865,1,L_SIZE),
				to_sfixed(0.9865,1,L_SIZE),
				to_sfixed(0.9865,1,L_SIZE),
				to_sfixed(0.9865,1,L_SIZE),
				to_sfixed(0.9865,1,L_SIZE),
				to_sfixed(0.9866,1,L_SIZE),
				to_sfixed(0.9866,1,L_SIZE),
				to_sfixed(0.9866,1,L_SIZE),
				to_sfixed(0.9866,1,L_SIZE),
				to_sfixed(0.9866,1,L_SIZE),
				to_sfixed(0.9866,1,L_SIZE),
				to_sfixed(0.9866,1,L_SIZE),
				to_sfixed(0.9866,1,L_SIZE),
				to_sfixed(0.9866,1,L_SIZE),
				to_sfixed(0.9866,1,L_SIZE),
				to_sfixed(0.9867,1,L_SIZE),
				to_sfixed(0.9867,1,L_SIZE),
				to_sfixed(0.9867,1,L_SIZE),
				to_sfixed(0.9867,1,L_SIZE),
				to_sfixed(0.9867,1,L_SIZE),
				to_sfixed(0.9867,1,L_SIZE),
				to_sfixed(0.9867,1,L_SIZE),
				to_sfixed(0.9867,1,L_SIZE),
				to_sfixed(0.9867,1,L_SIZE),
				to_sfixed(0.9867,1,L_SIZE),
				to_sfixed(0.9868,1,L_SIZE),
				to_sfixed(0.9868,1,L_SIZE),
				to_sfixed(0.9868,1,L_SIZE),
				to_sfixed(0.9868,1,L_SIZE),
				to_sfixed(0.9868,1,L_SIZE),
				to_sfixed(0.9868,1,L_SIZE),
				to_sfixed(0.9868,1,L_SIZE),
				to_sfixed(0.9868,1,L_SIZE),
				to_sfixed(0.9868,1,L_SIZE),
				to_sfixed(0.9868,1,L_SIZE),
				to_sfixed(0.9868,1,L_SIZE),
				to_sfixed(0.9869,1,L_SIZE),
				to_sfixed(0.9869,1,L_SIZE),
				to_sfixed(0.9869,1,L_SIZE),
				to_sfixed(0.9869,1,L_SIZE),
				to_sfixed(0.9869,1,L_SIZE),
				to_sfixed(0.9869,1,L_SIZE),
				to_sfixed(0.9869,1,L_SIZE),
				to_sfixed(0.9869,1,L_SIZE),
				to_sfixed(0.9869,1,L_SIZE),
				to_sfixed(0.9869,1,L_SIZE),
				to_sfixed(0.9870,1,L_SIZE),
				to_sfixed(0.9870,1,L_SIZE),
				to_sfixed(0.9870,1,L_SIZE),
				to_sfixed(0.9870,1,L_SIZE),
				to_sfixed(0.9870,1,L_SIZE),
				to_sfixed(0.9870,1,L_SIZE),
				to_sfixed(0.9870,1,L_SIZE),
				to_sfixed(0.9870,1,L_SIZE),
				to_sfixed(0.9870,1,L_SIZE),
				to_sfixed(0.9870,1,L_SIZE),
				to_sfixed(0.9870,1,L_SIZE),
				to_sfixed(0.9871,1,L_SIZE),
				to_sfixed(0.9871,1,L_SIZE),
				to_sfixed(0.9871,1,L_SIZE),
				to_sfixed(0.9871,1,L_SIZE),
				to_sfixed(0.9871,1,L_SIZE),
				to_sfixed(0.9871,1,L_SIZE),
				to_sfixed(0.9871,1,L_SIZE),
				to_sfixed(0.9871,1,L_SIZE),
				to_sfixed(0.9871,1,L_SIZE),
				to_sfixed(0.9871,1,L_SIZE),
				to_sfixed(0.9872,1,L_SIZE),
				to_sfixed(0.9872,1,L_SIZE),
				to_sfixed(0.9872,1,L_SIZE),
				to_sfixed(0.9872,1,L_SIZE),
				to_sfixed(0.9872,1,L_SIZE),
				to_sfixed(0.9872,1,L_SIZE),
				to_sfixed(0.9872,1,L_SIZE),
				to_sfixed(0.9872,1,L_SIZE),
				to_sfixed(0.9872,1,L_SIZE),
				to_sfixed(0.9872,1,L_SIZE),
				to_sfixed(0.9872,1,L_SIZE),
				to_sfixed(0.9873,1,L_SIZE),
				to_sfixed(0.9873,1,L_SIZE),
				to_sfixed(0.9873,1,L_SIZE),
				to_sfixed(0.9873,1,L_SIZE),
				to_sfixed(0.9873,1,L_SIZE),
				to_sfixed(0.9873,1,L_SIZE),
				to_sfixed(0.9873,1,L_SIZE),
				to_sfixed(0.9873,1,L_SIZE),
				to_sfixed(0.9873,1,L_SIZE),
				to_sfixed(0.9873,1,L_SIZE),
				to_sfixed(0.9873,1,L_SIZE),
				to_sfixed(0.9874,1,L_SIZE),
				to_sfixed(0.9874,1,L_SIZE),
				to_sfixed(0.9874,1,L_SIZE),
				to_sfixed(0.9874,1,L_SIZE),
				to_sfixed(0.9874,1,L_SIZE),
				to_sfixed(0.9874,1,L_SIZE),
				to_sfixed(0.9874,1,L_SIZE),
				to_sfixed(0.9874,1,L_SIZE),
				to_sfixed(0.9874,1,L_SIZE),
				to_sfixed(0.9874,1,L_SIZE),
				to_sfixed(0.9874,1,L_SIZE),
				to_sfixed(0.9875,1,L_SIZE),
				to_sfixed(0.9875,1,L_SIZE),
				to_sfixed(0.9875,1,L_SIZE),
				to_sfixed(0.9875,1,L_SIZE),
				to_sfixed(0.9875,1,L_SIZE),
				to_sfixed(0.9875,1,L_SIZE),
				to_sfixed(0.9875,1,L_SIZE),
				to_sfixed(0.9875,1,L_SIZE),
				to_sfixed(0.9875,1,L_SIZE),
				to_sfixed(0.9875,1,L_SIZE),
				to_sfixed(0.9875,1,L_SIZE),
				to_sfixed(0.9876,1,L_SIZE),
				to_sfixed(0.9876,1,L_SIZE),
				to_sfixed(0.9876,1,L_SIZE),
				to_sfixed(0.9876,1,L_SIZE),
				to_sfixed(0.9876,1,L_SIZE),
				to_sfixed(0.9876,1,L_SIZE),
				to_sfixed(0.9876,1,L_SIZE),
				to_sfixed(0.9876,1,L_SIZE),
				to_sfixed(0.9876,1,L_SIZE),
				to_sfixed(0.9876,1,L_SIZE),
				to_sfixed(0.9876,1,L_SIZE),
				to_sfixed(0.9877,1,L_SIZE),
				to_sfixed(0.9877,1,L_SIZE),
				to_sfixed(0.9877,1,L_SIZE),
				to_sfixed(0.9877,1,L_SIZE),
				to_sfixed(0.9877,1,L_SIZE),
				to_sfixed(0.9877,1,L_SIZE),
				to_sfixed(0.9877,1,L_SIZE),
				to_sfixed(0.9877,1,L_SIZE),
				to_sfixed(0.9877,1,L_SIZE),
				to_sfixed(0.9877,1,L_SIZE),
				to_sfixed(0.9877,1,L_SIZE),
				to_sfixed(0.9878,1,L_SIZE),
				to_sfixed(0.9878,1,L_SIZE),
				to_sfixed(0.9878,1,L_SIZE),
				to_sfixed(0.9878,1,L_SIZE),
				to_sfixed(0.9878,1,L_SIZE),
				to_sfixed(0.9878,1,L_SIZE),
				to_sfixed(0.9878,1,L_SIZE),
				to_sfixed(0.9878,1,L_SIZE),
				to_sfixed(0.9878,1,L_SIZE),
				to_sfixed(0.9878,1,L_SIZE),
				to_sfixed(0.9878,1,L_SIZE),
				to_sfixed(0.9879,1,L_SIZE),
				to_sfixed(0.9879,1,L_SIZE),
				to_sfixed(0.9879,1,L_SIZE),
				to_sfixed(0.9879,1,L_SIZE),
				to_sfixed(0.9879,1,L_SIZE),
				to_sfixed(0.9879,1,L_SIZE),
				to_sfixed(0.9879,1,L_SIZE),
				to_sfixed(0.9879,1,L_SIZE),
				to_sfixed(0.9879,1,L_SIZE),
				to_sfixed(0.9879,1,L_SIZE),
				to_sfixed(0.9879,1,L_SIZE),
				to_sfixed(0.9879,1,L_SIZE),
				to_sfixed(0.9880,1,L_SIZE),
				to_sfixed(0.9880,1,L_SIZE),
				to_sfixed(0.9880,1,L_SIZE),
				to_sfixed(0.9880,1,L_SIZE),
				to_sfixed(0.9880,1,L_SIZE),
				to_sfixed(0.9880,1,L_SIZE),
				to_sfixed(0.9880,1,L_SIZE),
				to_sfixed(0.9880,1,L_SIZE),
				to_sfixed(0.9880,1,L_SIZE),
				to_sfixed(0.9880,1,L_SIZE),
				to_sfixed(0.9880,1,L_SIZE),
				to_sfixed(0.9881,1,L_SIZE),
				to_sfixed(0.9881,1,L_SIZE),
				to_sfixed(0.9881,1,L_SIZE),
				to_sfixed(0.9881,1,L_SIZE),
				to_sfixed(0.9881,1,L_SIZE),
				to_sfixed(0.9881,1,L_SIZE),
				to_sfixed(0.9881,1,L_SIZE),
				to_sfixed(0.9881,1,L_SIZE),
				to_sfixed(0.9881,1,L_SIZE),
				to_sfixed(0.9881,1,L_SIZE),
				to_sfixed(0.9881,1,L_SIZE),
				to_sfixed(0.9881,1,L_SIZE),
				to_sfixed(0.9882,1,L_SIZE),
				to_sfixed(0.9882,1,L_SIZE),
				to_sfixed(0.9882,1,L_SIZE),
				to_sfixed(0.9882,1,L_SIZE),
				to_sfixed(0.9882,1,L_SIZE),
				to_sfixed(0.9882,1,L_SIZE),
				to_sfixed(0.9882,1,L_SIZE),
				to_sfixed(0.9882,1,L_SIZE),
				to_sfixed(0.9882,1,L_SIZE),
				to_sfixed(0.9882,1,L_SIZE),
				to_sfixed(0.9882,1,L_SIZE),
				to_sfixed(0.9883,1,L_SIZE),
				to_sfixed(0.9883,1,L_SIZE),
				to_sfixed(0.9883,1,L_SIZE),
				to_sfixed(0.9883,1,L_SIZE),
				to_sfixed(0.9883,1,L_SIZE),
				to_sfixed(0.9883,1,L_SIZE),
				to_sfixed(0.9883,1,L_SIZE),
				to_sfixed(0.9883,1,L_SIZE),
				to_sfixed(0.9883,1,L_SIZE),
				to_sfixed(0.9883,1,L_SIZE),
				to_sfixed(0.9883,1,L_SIZE),
				to_sfixed(0.9883,1,L_SIZE),
				to_sfixed(0.9884,1,L_SIZE),
				to_sfixed(0.9884,1,L_SIZE),
				to_sfixed(0.9884,1,L_SIZE),
				to_sfixed(0.9884,1,L_SIZE),
				to_sfixed(0.9884,1,L_SIZE),
				to_sfixed(0.9884,1,L_SIZE),
				to_sfixed(0.9884,1,L_SIZE),
				to_sfixed(0.9884,1,L_SIZE),
				to_sfixed(0.9884,1,L_SIZE),
				to_sfixed(0.9884,1,L_SIZE),
				to_sfixed(0.9884,1,L_SIZE),
				to_sfixed(0.9884,1,L_SIZE),
				to_sfixed(0.9885,1,L_SIZE),
				to_sfixed(0.9885,1,L_SIZE),
				to_sfixed(0.9885,1,L_SIZE),
				to_sfixed(0.9885,1,L_SIZE),
				to_sfixed(0.9885,1,L_SIZE),
				to_sfixed(0.9885,1,L_SIZE),
				to_sfixed(0.9885,1,L_SIZE),
				to_sfixed(0.9885,1,L_SIZE),
				to_sfixed(0.9885,1,L_SIZE),
				to_sfixed(0.9885,1,L_SIZE),
				to_sfixed(0.9885,1,L_SIZE),
				to_sfixed(0.9885,1,L_SIZE),
				to_sfixed(0.9886,1,L_SIZE),
				to_sfixed(0.9886,1,L_SIZE),
				to_sfixed(0.9886,1,L_SIZE),
				to_sfixed(0.9886,1,L_SIZE),
				to_sfixed(0.9886,1,L_SIZE),
				to_sfixed(0.9886,1,L_SIZE),
				to_sfixed(0.9886,1,L_SIZE),
				to_sfixed(0.9886,1,L_SIZE),
				to_sfixed(0.9886,1,L_SIZE),
				to_sfixed(0.9886,1,L_SIZE),
				to_sfixed(0.9886,1,L_SIZE),
				to_sfixed(0.9886,1,L_SIZE),
				to_sfixed(0.9887,1,L_SIZE),
				to_sfixed(0.9887,1,L_SIZE),
				to_sfixed(0.9887,1,L_SIZE),
				to_sfixed(0.9887,1,L_SIZE),
				to_sfixed(0.9887,1,L_SIZE),
				to_sfixed(0.9887,1,L_SIZE),
				to_sfixed(0.9887,1,L_SIZE),
				to_sfixed(0.9887,1,L_SIZE),
				to_sfixed(0.9887,1,L_SIZE),
				to_sfixed(0.9887,1,L_SIZE),
				to_sfixed(0.9887,1,L_SIZE),
				to_sfixed(0.9887,1,L_SIZE),
				to_sfixed(0.9888,1,L_SIZE),
				to_sfixed(0.9888,1,L_SIZE),
				to_sfixed(0.9888,1,L_SIZE),
				to_sfixed(0.9888,1,L_SIZE),
				to_sfixed(0.9888,1,L_SIZE),
				to_sfixed(0.9888,1,L_SIZE),
				to_sfixed(0.9888,1,L_SIZE),
				to_sfixed(0.9888,1,L_SIZE),
				to_sfixed(0.9888,1,L_SIZE),
				to_sfixed(0.9888,1,L_SIZE),
				to_sfixed(0.9888,1,L_SIZE),
				to_sfixed(0.9888,1,L_SIZE),
				to_sfixed(0.9889,1,L_SIZE),
				to_sfixed(0.9889,1,L_SIZE),
				to_sfixed(0.9889,1,L_SIZE),
				to_sfixed(0.9889,1,L_SIZE),
				to_sfixed(0.9889,1,L_SIZE),
				to_sfixed(0.9889,1,L_SIZE),
				to_sfixed(0.9889,1,L_SIZE),
				to_sfixed(0.9889,1,L_SIZE),
				to_sfixed(0.9889,1,L_SIZE),
				to_sfixed(0.9889,1,L_SIZE),
				to_sfixed(0.9889,1,L_SIZE),
				to_sfixed(0.9889,1,L_SIZE),
				to_sfixed(0.9889,1,L_SIZE),
				to_sfixed(0.9890,1,L_SIZE),
				to_sfixed(0.9890,1,L_SIZE),
				to_sfixed(0.9890,1,L_SIZE),
				to_sfixed(0.9890,1,L_SIZE),
				to_sfixed(0.9890,1,L_SIZE),
				to_sfixed(0.9890,1,L_SIZE),
				to_sfixed(0.9890,1,L_SIZE),
				to_sfixed(0.9890,1,L_SIZE),
				to_sfixed(0.9890,1,L_SIZE),
				to_sfixed(0.9890,1,L_SIZE),
				to_sfixed(0.9890,1,L_SIZE),
				to_sfixed(0.9890,1,L_SIZE),
				to_sfixed(0.9891,1,L_SIZE),
				to_sfixed(0.9891,1,L_SIZE),
				to_sfixed(0.9891,1,L_SIZE),
				to_sfixed(0.9891,1,L_SIZE),
				to_sfixed(0.9891,1,L_SIZE),
				to_sfixed(0.9891,1,L_SIZE),
				to_sfixed(0.9891,1,L_SIZE),
				to_sfixed(0.9891,1,L_SIZE),
				to_sfixed(0.9891,1,L_SIZE),
				to_sfixed(0.9891,1,L_SIZE),
				to_sfixed(0.9891,1,L_SIZE),
				to_sfixed(0.9891,1,L_SIZE),
				to_sfixed(0.9891,1,L_SIZE),
				to_sfixed(0.9892,1,L_SIZE),
				to_sfixed(0.9892,1,L_SIZE),
				to_sfixed(0.9892,1,L_SIZE),
				to_sfixed(0.9892,1,L_SIZE),
				to_sfixed(0.9892,1,L_SIZE),
				to_sfixed(0.9892,1,L_SIZE),
				to_sfixed(0.9892,1,L_SIZE),
				to_sfixed(0.9892,1,L_SIZE),
				to_sfixed(0.9892,1,L_SIZE),
				to_sfixed(0.9892,1,L_SIZE),
				to_sfixed(0.9892,1,L_SIZE),
				to_sfixed(0.9892,1,L_SIZE),
				to_sfixed(0.9893,1,L_SIZE),
				to_sfixed(0.9893,1,L_SIZE),
				to_sfixed(0.9893,1,L_SIZE),
				to_sfixed(0.9893,1,L_SIZE),
				to_sfixed(0.9893,1,L_SIZE),
				to_sfixed(0.9893,1,L_SIZE),
				to_sfixed(0.9893,1,L_SIZE),
				to_sfixed(0.9893,1,L_SIZE),
				to_sfixed(0.9893,1,L_SIZE),
				to_sfixed(0.9893,1,L_SIZE),
				to_sfixed(0.9893,1,L_SIZE),
				to_sfixed(0.9893,1,L_SIZE),
				to_sfixed(0.9893,1,L_SIZE),
				to_sfixed(0.9894,1,L_SIZE),
				to_sfixed(0.9894,1,L_SIZE),
				to_sfixed(0.9894,1,L_SIZE),
				to_sfixed(0.9894,1,L_SIZE),
				to_sfixed(0.9894,1,L_SIZE),
				to_sfixed(0.9894,1,L_SIZE),
				to_sfixed(0.9894,1,L_SIZE),
				to_sfixed(0.9894,1,L_SIZE),
				to_sfixed(0.9894,1,L_SIZE),
				to_sfixed(0.9894,1,L_SIZE),
				to_sfixed(0.9894,1,L_SIZE),
				to_sfixed(0.9894,1,L_SIZE),
				to_sfixed(0.9894,1,L_SIZE),
				to_sfixed(0.9895,1,L_SIZE),
				to_sfixed(0.9895,1,L_SIZE),
				to_sfixed(0.9895,1,L_SIZE),
				to_sfixed(0.9895,1,L_SIZE),
				to_sfixed(0.9895,1,L_SIZE),
				to_sfixed(0.9895,1,L_SIZE),
				to_sfixed(0.9895,1,L_SIZE),
				to_sfixed(0.9895,1,L_SIZE),
				to_sfixed(0.9895,1,L_SIZE),
				to_sfixed(0.9895,1,L_SIZE),
				to_sfixed(0.9895,1,L_SIZE),
				to_sfixed(0.9895,1,L_SIZE),
				to_sfixed(0.9895,1,L_SIZE),
				to_sfixed(0.9896,1,L_SIZE),
				to_sfixed(0.9896,1,L_SIZE),
				to_sfixed(0.9896,1,L_SIZE),
				to_sfixed(0.9896,1,L_SIZE),
				to_sfixed(0.9896,1,L_SIZE),
				to_sfixed(0.9896,1,L_SIZE),
				to_sfixed(0.9896,1,L_SIZE),
				to_sfixed(0.9896,1,L_SIZE),
				to_sfixed(0.9896,1,L_SIZE),
				to_sfixed(0.9896,1,L_SIZE),
				to_sfixed(0.9896,1,L_SIZE),
				to_sfixed(0.9896,1,L_SIZE),
				to_sfixed(0.9896,1,L_SIZE),
				to_sfixed(0.9897,1,L_SIZE),
				to_sfixed(0.9897,1,L_SIZE),
				to_sfixed(0.9897,1,L_SIZE),
				to_sfixed(0.9897,1,L_SIZE),
				to_sfixed(0.9897,1,L_SIZE),
				to_sfixed(0.9897,1,L_SIZE),
				to_sfixed(0.9897,1,L_SIZE),
				to_sfixed(0.9897,1,L_SIZE),
				to_sfixed(0.9897,1,L_SIZE),
				to_sfixed(0.9897,1,L_SIZE),
				to_sfixed(0.9897,1,L_SIZE),
				to_sfixed(0.9897,1,L_SIZE),
				to_sfixed(0.9897,1,L_SIZE),
				to_sfixed(0.9897,1,L_SIZE),
				to_sfixed(0.9898,1,L_SIZE),
				to_sfixed(0.9898,1,L_SIZE),
				to_sfixed(0.9898,1,L_SIZE),
				to_sfixed(0.9898,1,L_SIZE),
				to_sfixed(0.9898,1,L_SIZE),
				to_sfixed(0.9898,1,L_SIZE),
				to_sfixed(0.9898,1,L_SIZE),
				to_sfixed(0.9898,1,L_SIZE),
				to_sfixed(0.9898,1,L_SIZE),
				to_sfixed(0.9898,1,L_SIZE),
				to_sfixed(0.9898,1,L_SIZE),
				to_sfixed(0.9898,1,L_SIZE),
				to_sfixed(0.9898,1,L_SIZE),
				to_sfixed(0.9899,1,L_SIZE),
				to_sfixed(0.9899,1,L_SIZE),
				to_sfixed(0.9899,1,L_SIZE),
				to_sfixed(0.9899,1,L_SIZE),
				to_sfixed(0.9899,1,L_SIZE),
				to_sfixed(0.9899,1,L_SIZE),
				to_sfixed(0.9899,1,L_SIZE),
				to_sfixed(0.9899,1,L_SIZE),
				to_sfixed(0.9899,1,L_SIZE),
				to_sfixed(0.9899,1,L_SIZE),
				to_sfixed(0.9899,1,L_SIZE),
				to_sfixed(0.9899,1,L_SIZE),
				to_sfixed(0.9899,1,L_SIZE),
				to_sfixed(0.9899,1,L_SIZE),
				to_sfixed(0.9900,1,L_SIZE),
				to_sfixed(0.9900,1,L_SIZE),
				to_sfixed(0.9900,1,L_SIZE),
				to_sfixed(0.9900,1,L_SIZE),
				to_sfixed(0.9900,1,L_SIZE),
				to_sfixed(0.9900,1,L_SIZE),
				to_sfixed(0.9900,1,L_SIZE),
				to_sfixed(0.9900,1,L_SIZE),
				to_sfixed(0.9900,1,L_SIZE),
				to_sfixed(0.9900,1,L_SIZE),
				to_sfixed(0.9900,1,L_SIZE),
				to_sfixed(0.9900,1,L_SIZE),
				to_sfixed(0.9900,1,L_SIZE),
				to_sfixed(0.9900,1,L_SIZE),
				to_sfixed(0.9901,1,L_SIZE),
				to_sfixed(0.9901,1,L_SIZE),
				to_sfixed(0.9901,1,L_SIZE),
				to_sfixed(0.9901,1,L_SIZE),
				to_sfixed(0.9901,1,L_SIZE),
				to_sfixed(0.9901,1,L_SIZE),
				to_sfixed(0.9901,1,L_SIZE),
				to_sfixed(0.9901,1,L_SIZE),
				to_sfixed(0.9901,1,L_SIZE),
				to_sfixed(0.9901,1,L_SIZE),
				to_sfixed(0.9901,1,L_SIZE),
				to_sfixed(0.9901,1,L_SIZE),
				to_sfixed(0.9901,1,L_SIZE),
				to_sfixed(0.9902,1,L_SIZE),
				to_sfixed(0.9902,1,L_SIZE),
				to_sfixed(0.9902,1,L_SIZE),
				to_sfixed(0.9902,1,L_SIZE),
				to_sfixed(0.9902,1,L_SIZE),
				to_sfixed(0.9902,1,L_SIZE),
				to_sfixed(0.9902,1,L_SIZE),
				to_sfixed(0.9902,1,L_SIZE),
				to_sfixed(0.9902,1,L_SIZE),
				to_sfixed(0.9902,1,L_SIZE),
				to_sfixed(0.9902,1,L_SIZE),
				to_sfixed(0.9902,1,L_SIZE),
				to_sfixed(0.9902,1,L_SIZE),
				to_sfixed(0.9902,1,L_SIZE),
				to_sfixed(0.9903,1,L_SIZE),
				to_sfixed(0.9903,1,L_SIZE),
				to_sfixed(0.9903,1,L_SIZE),
				to_sfixed(0.9903,1,L_SIZE),
				to_sfixed(0.9903,1,L_SIZE),
				to_sfixed(0.9903,1,L_SIZE),
				to_sfixed(0.9903,1,L_SIZE),
				to_sfixed(0.9903,1,L_SIZE),
				to_sfixed(0.9903,1,L_SIZE),
				to_sfixed(0.9903,1,L_SIZE),
				to_sfixed(0.9903,1,L_SIZE),
				to_sfixed(0.9903,1,L_SIZE),
				to_sfixed(0.9903,1,L_SIZE),
				to_sfixed(0.9903,1,L_SIZE),
				to_sfixed(0.9903,1,L_SIZE),
				to_sfixed(0.9904,1,L_SIZE),
				to_sfixed(0.9904,1,L_SIZE),
				to_sfixed(0.9904,1,L_SIZE),
				to_sfixed(0.9904,1,L_SIZE),
				to_sfixed(0.9904,1,L_SIZE),
				to_sfixed(0.9904,1,L_SIZE),
				to_sfixed(0.9904,1,L_SIZE),
				to_sfixed(0.9904,1,L_SIZE),
				to_sfixed(0.9904,1,L_SIZE),
				to_sfixed(0.9904,1,L_SIZE),
				to_sfixed(0.9904,1,L_SIZE),
				to_sfixed(0.9904,1,L_SIZE),
				to_sfixed(0.9904,1,L_SIZE),
				to_sfixed(0.9904,1,L_SIZE),
				to_sfixed(0.9905,1,L_SIZE),
				to_sfixed(0.9905,1,L_SIZE),
				to_sfixed(0.9905,1,L_SIZE),
				to_sfixed(0.9905,1,L_SIZE),
				to_sfixed(0.9905,1,L_SIZE),
				to_sfixed(0.9905,1,L_SIZE),
				to_sfixed(0.9905,1,L_SIZE),
				to_sfixed(0.9905,1,L_SIZE),
				to_sfixed(0.9905,1,L_SIZE),
				to_sfixed(0.9905,1,L_SIZE),
				to_sfixed(0.9905,1,L_SIZE),
				to_sfixed(0.9905,1,L_SIZE),
				to_sfixed(0.9905,1,L_SIZE),
				to_sfixed(0.9905,1,L_SIZE),
				to_sfixed(0.9906,1,L_SIZE),
				to_sfixed(0.9906,1,L_SIZE),
				to_sfixed(0.9906,1,L_SIZE),
				to_sfixed(0.9906,1,L_SIZE),
				to_sfixed(0.9906,1,L_SIZE),
				to_sfixed(0.9906,1,L_SIZE),
				to_sfixed(0.9906,1,L_SIZE),
				to_sfixed(0.9906,1,L_SIZE),
				to_sfixed(0.9906,1,L_SIZE),
				to_sfixed(0.9906,1,L_SIZE),
				to_sfixed(0.9906,1,L_SIZE),
				to_sfixed(0.9906,1,L_SIZE),
				to_sfixed(0.9906,1,L_SIZE),
				to_sfixed(0.9906,1,L_SIZE),
				to_sfixed(0.9906,1,L_SIZE),
				to_sfixed(0.9907,1,L_SIZE),
				to_sfixed(0.9907,1,L_SIZE),
				to_sfixed(0.9907,1,L_SIZE),
				to_sfixed(0.9907,1,L_SIZE),
				to_sfixed(0.9907,1,L_SIZE),
				to_sfixed(0.9907,1,L_SIZE),
				to_sfixed(0.9907,1,L_SIZE),
				to_sfixed(0.9907,1,L_SIZE),
				to_sfixed(0.9907,1,L_SIZE),
				to_sfixed(0.9907,1,L_SIZE),
				to_sfixed(0.9907,1,L_SIZE),
				to_sfixed(0.9907,1,L_SIZE),
				to_sfixed(0.9907,1,L_SIZE),
				to_sfixed(0.9907,1,L_SIZE),
				to_sfixed(0.9907,1,L_SIZE),
				to_sfixed(0.9908,1,L_SIZE),
				to_sfixed(0.9908,1,L_SIZE),
				to_sfixed(0.9908,1,L_SIZE),
				to_sfixed(0.9908,1,L_SIZE),
				to_sfixed(0.9908,1,L_SIZE),
				to_sfixed(0.9908,1,L_SIZE),
				to_sfixed(0.9908,1,L_SIZE),
				to_sfixed(0.9908,1,L_SIZE),
				to_sfixed(0.9908,1,L_SIZE),
				to_sfixed(0.9908,1,L_SIZE),
				to_sfixed(0.9908,1,L_SIZE),
				to_sfixed(0.9908,1,L_SIZE),
				to_sfixed(0.9908,1,L_SIZE),
				to_sfixed(0.9908,1,L_SIZE),
				to_sfixed(0.9909,1,L_SIZE),
				to_sfixed(0.9909,1,L_SIZE),
				to_sfixed(0.9909,1,L_SIZE),
				to_sfixed(0.9909,1,L_SIZE),
				to_sfixed(0.9909,1,L_SIZE),
				to_sfixed(0.9909,1,L_SIZE),
				to_sfixed(0.9909,1,L_SIZE),
				to_sfixed(0.9909,1,L_SIZE),
				to_sfixed(0.9909,1,L_SIZE),
				to_sfixed(0.9909,1,L_SIZE),
				to_sfixed(0.9909,1,L_SIZE),
				to_sfixed(0.9909,1,L_SIZE),
				to_sfixed(0.9909,1,L_SIZE),
				to_sfixed(0.9909,1,L_SIZE),
				to_sfixed(0.9909,1,L_SIZE),
				to_sfixed(0.9909,1,L_SIZE),
				to_sfixed(0.9910,1,L_SIZE),
				to_sfixed(0.9910,1,L_SIZE),
				to_sfixed(0.9910,1,L_SIZE),
				to_sfixed(0.9910,1,L_SIZE),
				to_sfixed(0.9910,1,L_SIZE),
				to_sfixed(0.9910,1,L_SIZE),
				to_sfixed(0.9910,1,L_SIZE),
				to_sfixed(0.9910,1,L_SIZE),
				to_sfixed(0.9910,1,L_SIZE),
				to_sfixed(0.9910,1,L_SIZE),
				to_sfixed(0.9910,1,L_SIZE),
				to_sfixed(0.9910,1,L_SIZE),
				to_sfixed(0.9910,1,L_SIZE),
				to_sfixed(0.9910,1,L_SIZE),
				to_sfixed(0.9910,1,L_SIZE),
				to_sfixed(0.9911,1,L_SIZE),
				to_sfixed(0.9911,1,L_SIZE),
				to_sfixed(0.9911,1,L_SIZE),
				to_sfixed(0.9911,1,L_SIZE),
				to_sfixed(0.9911,1,L_SIZE),
				to_sfixed(0.9911,1,L_SIZE),
				to_sfixed(0.9911,1,L_SIZE),
				to_sfixed(0.9911,1,L_SIZE),
				to_sfixed(0.9911,1,L_SIZE),
				to_sfixed(0.9911,1,L_SIZE),
				to_sfixed(0.9911,1,L_SIZE),
				to_sfixed(0.9911,1,L_SIZE),
				to_sfixed(0.9911,1,L_SIZE),
				to_sfixed(0.9911,1,L_SIZE),
				to_sfixed(0.9911,1,L_SIZE),
				to_sfixed(0.9912,1,L_SIZE),
				to_sfixed(0.9912,1,L_SIZE),
				to_sfixed(0.9912,1,L_SIZE),
				to_sfixed(0.9912,1,L_SIZE),
				to_sfixed(0.9912,1,L_SIZE),
				to_sfixed(0.9912,1,L_SIZE),
				to_sfixed(0.9912,1,L_SIZE),
				to_sfixed(0.9912,1,L_SIZE),
				to_sfixed(0.9912,1,L_SIZE),
				to_sfixed(0.9912,1,L_SIZE),
				to_sfixed(0.9912,1,L_SIZE),
				to_sfixed(0.9912,1,L_SIZE),
				to_sfixed(0.9912,1,L_SIZE),
				to_sfixed(0.9912,1,L_SIZE),
				to_sfixed(0.9912,1,L_SIZE),
				to_sfixed(0.9912,1,L_SIZE),
				to_sfixed(0.9913,1,L_SIZE),
				to_sfixed(0.9913,1,L_SIZE),
				to_sfixed(0.9913,1,L_SIZE),
				to_sfixed(0.9913,1,L_SIZE),
				to_sfixed(0.9913,1,L_SIZE),
				to_sfixed(0.9913,1,L_SIZE),
				to_sfixed(0.9913,1,L_SIZE),
				to_sfixed(0.9913,1,L_SIZE),
				to_sfixed(0.9913,1,L_SIZE),
				to_sfixed(0.9913,1,L_SIZE),
				to_sfixed(0.9913,1,L_SIZE),
				to_sfixed(0.9913,1,L_SIZE),
				to_sfixed(0.9913,1,L_SIZE),
				to_sfixed(0.9913,1,L_SIZE),
				to_sfixed(0.9913,1,L_SIZE),
				to_sfixed(0.9913,1,L_SIZE),
				to_sfixed(0.9914,1,L_SIZE),
				to_sfixed(0.9914,1,L_SIZE),
				to_sfixed(0.9914,1,L_SIZE),
				to_sfixed(0.9914,1,L_SIZE),
				to_sfixed(0.9914,1,L_SIZE),
				to_sfixed(0.9914,1,L_SIZE),
				to_sfixed(0.9914,1,L_SIZE),
				to_sfixed(0.9914,1,L_SIZE),
				to_sfixed(0.9914,1,L_SIZE),
				to_sfixed(0.9914,1,L_SIZE),
				to_sfixed(0.9914,1,L_SIZE),
				to_sfixed(0.9914,1,L_SIZE),
				to_sfixed(0.9914,1,L_SIZE),
				to_sfixed(0.9914,1,L_SIZE),
				to_sfixed(0.9914,1,L_SIZE),
				to_sfixed(0.9914,1,L_SIZE),
				to_sfixed(0.9915,1,L_SIZE),
				to_sfixed(0.9915,1,L_SIZE),
				to_sfixed(0.9915,1,L_SIZE),
				to_sfixed(0.9915,1,L_SIZE),
				to_sfixed(0.9915,1,L_SIZE),
				to_sfixed(0.9915,1,L_SIZE),
				to_sfixed(0.9915,1,L_SIZE),
				to_sfixed(0.9915,1,L_SIZE),
				to_sfixed(0.9915,1,L_SIZE),
				to_sfixed(0.9915,1,L_SIZE),
				to_sfixed(0.9915,1,L_SIZE),
				to_sfixed(0.9915,1,L_SIZE),
				to_sfixed(0.9915,1,L_SIZE),
				to_sfixed(0.9915,1,L_SIZE),
				to_sfixed(0.9915,1,L_SIZE),
				to_sfixed(0.9915,1,L_SIZE),
				to_sfixed(0.9916,1,L_SIZE),
				to_sfixed(0.9916,1,L_SIZE),
				to_sfixed(0.9916,1,L_SIZE),
				to_sfixed(0.9916,1,L_SIZE),
				to_sfixed(0.9916,1,L_SIZE),
				to_sfixed(0.9916,1,L_SIZE),
				to_sfixed(0.9916,1,L_SIZE),
				to_sfixed(0.9916,1,L_SIZE),
				to_sfixed(0.9916,1,L_SIZE),
				to_sfixed(0.9916,1,L_SIZE),
				to_sfixed(0.9916,1,L_SIZE),
				to_sfixed(0.9916,1,L_SIZE),
				to_sfixed(0.9916,1,L_SIZE),
				to_sfixed(0.9916,1,L_SIZE),
				to_sfixed(0.9916,1,L_SIZE),
				to_sfixed(0.9916,1,L_SIZE),
				to_sfixed(0.9917,1,L_SIZE),
				to_sfixed(0.9917,1,L_SIZE),
				to_sfixed(0.9917,1,L_SIZE),
				to_sfixed(0.9917,1,L_SIZE),
				to_sfixed(0.9917,1,L_SIZE),
				to_sfixed(0.9917,1,L_SIZE),
				to_sfixed(0.9917,1,L_SIZE),
				to_sfixed(0.9917,1,L_SIZE),
				to_sfixed(0.9917,1,L_SIZE),
				to_sfixed(0.9917,1,L_SIZE),
				to_sfixed(0.9917,1,L_SIZE),
				to_sfixed(0.9917,1,L_SIZE),
				to_sfixed(0.9917,1,L_SIZE),
				to_sfixed(0.9917,1,L_SIZE),
				to_sfixed(0.9917,1,L_SIZE),
				to_sfixed(0.9917,1,L_SIZE),
				to_sfixed(0.9918,1,L_SIZE),
				to_sfixed(0.9918,1,L_SIZE),
				to_sfixed(0.9918,1,L_SIZE),
				to_sfixed(0.9918,1,L_SIZE),
				to_sfixed(0.9918,1,L_SIZE),
				to_sfixed(0.9918,1,L_SIZE),
				to_sfixed(0.9918,1,L_SIZE),
				to_sfixed(0.9918,1,L_SIZE),
				to_sfixed(0.9918,1,L_SIZE),
				to_sfixed(0.9918,1,L_SIZE),
				to_sfixed(0.9918,1,L_SIZE),
				to_sfixed(0.9918,1,L_SIZE),
				to_sfixed(0.9918,1,L_SIZE),
				to_sfixed(0.9918,1,L_SIZE),
				to_sfixed(0.9918,1,L_SIZE),
				to_sfixed(0.9918,1,L_SIZE),
				to_sfixed(0.9918,1,L_SIZE),
				to_sfixed(0.9919,1,L_SIZE),
				to_sfixed(0.9919,1,L_SIZE),
				to_sfixed(0.9919,1,L_SIZE),
				to_sfixed(0.9919,1,L_SIZE),
				to_sfixed(0.9919,1,L_SIZE),
				to_sfixed(0.9919,1,L_SIZE),
				to_sfixed(0.9919,1,L_SIZE),
				to_sfixed(0.9919,1,L_SIZE),
				to_sfixed(0.9919,1,L_SIZE),
				to_sfixed(0.9919,1,L_SIZE),
				to_sfixed(0.9919,1,L_SIZE),
				to_sfixed(0.9919,1,L_SIZE),
				to_sfixed(0.9919,1,L_SIZE),
				to_sfixed(0.9919,1,L_SIZE),
				to_sfixed(0.9919,1,L_SIZE),
				to_sfixed(0.9919,1,L_SIZE),
				to_sfixed(0.9919,1,L_SIZE),
				to_sfixed(0.9920,1,L_SIZE),
				to_sfixed(0.9920,1,L_SIZE),
				to_sfixed(0.9920,1,L_SIZE),
				to_sfixed(0.9920,1,L_SIZE),
				to_sfixed(0.9920,1,L_SIZE),
				to_sfixed(0.9920,1,L_SIZE),
				to_sfixed(0.9920,1,L_SIZE),
				to_sfixed(0.9920,1,L_SIZE),
				to_sfixed(0.9920,1,L_SIZE),
				to_sfixed(0.9920,1,L_SIZE),
				to_sfixed(0.9920,1,L_SIZE),
				to_sfixed(0.9920,1,L_SIZE),
				to_sfixed(0.9920,1,L_SIZE),
				to_sfixed(0.9920,1,L_SIZE),
				to_sfixed(0.9920,1,L_SIZE),
				to_sfixed(0.9920,1,L_SIZE),
				to_sfixed(0.9920,1,L_SIZE),
				to_sfixed(0.9921,1,L_SIZE),
				to_sfixed(0.9921,1,L_SIZE),
				to_sfixed(0.9921,1,L_SIZE),
				to_sfixed(0.9921,1,L_SIZE),
				to_sfixed(0.9921,1,L_SIZE),
				to_sfixed(0.9921,1,L_SIZE),
				to_sfixed(0.9921,1,L_SIZE),
				to_sfixed(0.9921,1,L_SIZE),
				to_sfixed(0.9921,1,L_SIZE),
				to_sfixed(0.9921,1,L_SIZE),
				to_sfixed(0.9921,1,L_SIZE),
				to_sfixed(0.9921,1,L_SIZE),
				to_sfixed(0.9921,1,L_SIZE),
				to_sfixed(0.9921,1,L_SIZE),
				to_sfixed(0.9921,1,L_SIZE),
				to_sfixed(0.9921,1,L_SIZE),
				to_sfixed(0.9921,1,L_SIZE),
				to_sfixed(0.9921,1,L_SIZE),
				to_sfixed(0.9922,1,L_SIZE),
				to_sfixed(0.9922,1,L_SIZE),
				to_sfixed(0.9922,1,L_SIZE),
				to_sfixed(0.9922,1,L_SIZE),
				to_sfixed(0.9922,1,L_SIZE),
				to_sfixed(0.9922,1,L_SIZE),
				to_sfixed(0.9922,1,L_SIZE),
				to_sfixed(0.9922,1,L_SIZE),
				to_sfixed(0.9922,1,L_SIZE),
				to_sfixed(0.9922,1,L_SIZE),
				to_sfixed(0.9922,1,L_SIZE),
				to_sfixed(0.9922,1,L_SIZE),
				to_sfixed(0.9922,1,L_SIZE),
				to_sfixed(0.9922,1,L_SIZE),
				to_sfixed(0.9922,1,L_SIZE),
				to_sfixed(0.9922,1,L_SIZE),
				to_sfixed(0.9922,1,L_SIZE),
				to_sfixed(0.9923,1,L_SIZE),
				to_sfixed(0.9923,1,L_SIZE),
				to_sfixed(0.9923,1,L_SIZE),
				to_sfixed(0.9923,1,L_SIZE),
				to_sfixed(0.9923,1,L_SIZE),
				to_sfixed(0.9923,1,L_SIZE),
				to_sfixed(0.9923,1,L_SIZE),
				to_sfixed(0.9923,1,L_SIZE),
				to_sfixed(0.9923,1,L_SIZE),
				to_sfixed(0.9923,1,L_SIZE),
				to_sfixed(0.9923,1,L_SIZE),
				to_sfixed(0.9923,1,L_SIZE),
				to_sfixed(0.9923,1,L_SIZE),
				to_sfixed(0.9923,1,L_SIZE),
				to_sfixed(0.9923,1,L_SIZE),
				to_sfixed(0.9923,1,L_SIZE),
				to_sfixed(0.9923,1,L_SIZE),
				to_sfixed(0.9923,1,L_SIZE),
				to_sfixed(0.9924,1,L_SIZE),
				to_sfixed(0.9924,1,L_SIZE),
				to_sfixed(0.9924,1,L_SIZE),
				to_sfixed(0.9924,1,L_SIZE),
				to_sfixed(0.9924,1,L_SIZE),
				to_sfixed(0.9924,1,L_SIZE),
				to_sfixed(0.9924,1,L_SIZE),
				to_sfixed(0.9924,1,L_SIZE),
				to_sfixed(0.9924,1,L_SIZE),
				to_sfixed(0.9924,1,L_SIZE),
				to_sfixed(0.9924,1,L_SIZE),
				to_sfixed(0.9924,1,L_SIZE),
				to_sfixed(0.9924,1,L_SIZE),
				to_sfixed(0.9924,1,L_SIZE),
				to_sfixed(0.9924,1,L_SIZE),
				to_sfixed(0.9924,1,L_SIZE),
				to_sfixed(0.9924,1,L_SIZE),
				to_sfixed(0.9924,1,L_SIZE),
				to_sfixed(0.9925,1,L_SIZE),
				to_sfixed(0.9925,1,L_SIZE),
				to_sfixed(0.9925,1,L_SIZE),
				to_sfixed(0.9925,1,L_SIZE),
				to_sfixed(0.9925,1,L_SIZE),
				to_sfixed(0.9925,1,L_SIZE),
				to_sfixed(0.9925,1,L_SIZE),
				to_sfixed(0.9925,1,L_SIZE),
				to_sfixed(0.9925,1,L_SIZE),
				to_sfixed(0.9925,1,L_SIZE),
				to_sfixed(0.9925,1,L_SIZE),
				to_sfixed(0.9925,1,L_SIZE),
				to_sfixed(0.9925,1,L_SIZE),
				to_sfixed(0.9925,1,L_SIZE),
				to_sfixed(0.9925,1,L_SIZE),
				to_sfixed(0.9925,1,L_SIZE),
				to_sfixed(0.9925,1,L_SIZE),
				to_sfixed(0.9925,1,L_SIZE),
				to_sfixed(0.9926,1,L_SIZE),
				to_sfixed(0.9926,1,L_SIZE),
				to_sfixed(0.9926,1,L_SIZE),
				to_sfixed(0.9926,1,L_SIZE),
				to_sfixed(0.9926,1,L_SIZE),
				to_sfixed(0.9926,1,L_SIZE),
				to_sfixed(0.9926,1,L_SIZE),
				to_sfixed(0.9926,1,L_SIZE),
				to_sfixed(0.9926,1,L_SIZE),
				to_sfixed(0.9926,1,L_SIZE),
				to_sfixed(0.9926,1,L_SIZE),
				to_sfixed(0.9926,1,L_SIZE),
				to_sfixed(0.9926,1,L_SIZE),
				to_sfixed(0.9926,1,L_SIZE),
				to_sfixed(0.9926,1,L_SIZE),
				to_sfixed(0.9926,1,L_SIZE),
				to_sfixed(0.9926,1,L_SIZE),
				to_sfixed(0.9926,1,L_SIZE),
				to_sfixed(0.9926,1,L_SIZE),
				to_sfixed(0.9927,1,L_SIZE),
				to_sfixed(0.9927,1,L_SIZE),
				to_sfixed(0.9927,1,L_SIZE),
				to_sfixed(0.9927,1,L_SIZE),
				to_sfixed(0.9927,1,L_SIZE),
				to_sfixed(0.9927,1,L_SIZE),
				to_sfixed(0.9927,1,L_SIZE),
				to_sfixed(0.9927,1,L_SIZE),
				to_sfixed(0.9927,1,L_SIZE),
				to_sfixed(0.9927,1,L_SIZE),
				to_sfixed(0.9927,1,L_SIZE),
				to_sfixed(0.9927,1,L_SIZE),
				to_sfixed(0.9927,1,L_SIZE),
				to_sfixed(0.9927,1,L_SIZE),
				to_sfixed(0.9927,1,L_SIZE),
				to_sfixed(0.9927,1,L_SIZE),
				to_sfixed(0.9927,1,L_SIZE),
				to_sfixed(0.9927,1,L_SIZE),
				to_sfixed(0.9927,1,L_SIZE),
				to_sfixed(0.9928,1,L_SIZE),
				to_sfixed(0.9928,1,L_SIZE),
				to_sfixed(0.9928,1,L_SIZE),
				to_sfixed(0.9928,1,L_SIZE),
				to_sfixed(0.9928,1,L_SIZE),
				to_sfixed(0.9928,1,L_SIZE),
				to_sfixed(0.9928,1,L_SIZE),
				to_sfixed(0.9928,1,L_SIZE),
				to_sfixed(0.9928,1,L_SIZE),
				to_sfixed(0.9928,1,L_SIZE),
				to_sfixed(0.9928,1,L_SIZE),
				to_sfixed(0.9928,1,L_SIZE),
				to_sfixed(0.9928,1,L_SIZE),
				to_sfixed(0.9928,1,L_SIZE),
				to_sfixed(0.9928,1,L_SIZE),
				to_sfixed(0.9928,1,L_SIZE),
				to_sfixed(0.9928,1,L_SIZE),
				to_sfixed(0.9928,1,L_SIZE),
				to_sfixed(0.9928,1,L_SIZE),
				to_sfixed(0.9929,1,L_SIZE),
				to_sfixed(0.9929,1,L_SIZE),
				to_sfixed(0.9929,1,L_SIZE),
				to_sfixed(0.9929,1,L_SIZE),
				to_sfixed(0.9929,1,L_SIZE),
				to_sfixed(0.9929,1,L_SIZE),
				to_sfixed(0.9929,1,L_SIZE),
				to_sfixed(0.9929,1,L_SIZE),
				to_sfixed(0.9929,1,L_SIZE),
				to_sfixed(0.9929,1,L_SIZE),
				to_sfixed(0.9929,1,L_SIZE),
				to_sfixed(0.9929,1,L_SIZE),
				to_sfixed(0.9929,1,L_SIZE),
				to_sfixed(0.9929,1,L_SIZE),
				to_sfixed(0.9929,1,L_SIZE),
				to_sfixed(0.9929,1,L_SIZE),
				to_sfixed(0.9929,1,L_SIZE),
				to_sfixed(0.9929,1,L_SIZE),
				to_sfixed(0.9929,1,L_SIZE),
				to_sfixed(0.9930,1,L_SIZE),
				to_sfixed(0.9930,1,L_SIZE),
				to_sfixed(0.9930,1,L_SIZE),
				to_sfixed(0.9930,1,L_SIZE),
				to_sfixed(0.9930,1,L_SIZE),
				to_sfixed(0.9930,1,L_SIZE),
				to_sfixed(0.9930,1,L_SIZE),
				to_sfixed(0.9930,1,L_SIZE),
				to_sfixed(0.9930,1,L_SIZE),
				to_sfixed(0.9930,1,L_SIZE),
				to_sfixed(0.9930,1,L_SIZE),
				to_sfixed(0.9930,1,L_SIZE),
				to_sfixed(0.9930,1,L_SIZE),
				to_sfixed(0.9930,1,L_SIZE),
				to_sfixed(0.9930,1,L_SIZE),
				to_sfixed(0.9930,1,L_SIZE),
				to_sfixed(0.9930,1,L_SIZE),
				to_sfixed(0.9930,1,L_SIZE),
				to_sfixed(0.9930,1,L_SIZE),
				to_sfixed(0.9931,1,L_SIZE),
				to_sfixed(0.9931,1,L_SIZE),
				to_sfixed(0.9931,1,L_SIZE),
				to_sfixed(0.9931,1,L_SIZE),
				to_sfixed(0.9931,1,L_SIZE),
				to_sfixed(0.9931,1,L_SIZE),
				to_sfixed(0.9931,1,L_SIZE),
				to_sfixed(0.9931,1,L_SIZE),
				to_sfixed(0.9931,1,L_SIZE),
				to_sfixed(0.9931,1,L_SIZE),
				to_sfixed(0.9931,1,L_SIZE),
				to_sfixed(0.9931,1,L_SIZE),
				to_sfixed(0.9931,1,L_SIZE),
				to_sfixed(0.9931,1,L_SIZE),
				to_sfixed(0.9931,1,L_SIZE),
				to_sfixed(0.9931,1,L_SIZE),
				to_sfixed(0.9931,1,L_SIZE),
				to_sfixed(0.9931,1,L_SIZE),
				to_sfixed(0.9931,1,L_SIZE),
				to_sfixed(0.9931,1,L_SIZE),
				to_sfixed(0.9932,1,L_SIZE),
				to_sfixed(0.9932,1,L_SIZE),
				to_sfixed(0.9932,1,L_SIZE),
				to_sfixed(0.9932,1,L_SIZE),
				to_sfixed(0.9932,1,L_SIZE),
				to_sfixed(0.9932,1,L_SIZE),
				to_sfixed(0.9932,1,L_SIZE),
				to_sfixed(0.9932,1,L_SIZE),
				to_sfixed(0.9932,1,L_SIZE),
				to_sfixed(0.9932,1,L_SIZE),
				to_sfixed(0.9932,1,L_SIZE),
				to_sfixed(0.9932,1,L_SIZE),
				to_sfixed(0.9932,1,L_SIZE),
				to_sfixed(0.9932,1,L_SIZE),
				to_sfixed(0.9932,1,L_SIZE),
				to_sfixed(0.9932,1,L_SIZE),
				to_sfixed(0.9932,1,L_SIZE),
				to_sfixed(0.9932,1,L_SIZE),
				to_sfixed(0.9932,1,L_SIZE),
				to_sfixed(0.9932,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9933,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9934,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9935,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9936,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9937,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9938,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9939,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9940,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9941,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9942,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9943,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9944,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9945,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9946,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9947,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9948,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9949,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9950,1,L_SIZE),
				to_sfixed(0.9951,1,L_SIZE)
			);
	  -- Signals
	signal IN_UNSIGNED						: unsigned(13 downto 0);
	signal LOOKUP_TABLE_K 					: unsigned(13 downto 0);
	signal LOOKUP_TABLE_OUT 				: INPUT_SFIXED;
	signal LOOKUP_TABLE_OUT_CONSTRAINED	: CONSTRAINED_SFIXED;
	signal UNIT_DELAY_OUT					: CONSTRAINED_SFIXED;
	
	
--=============================================================================
-- architecture begin
--=============================================================================	
	begin
		IN_UNSIGNED <= unsigned(X_VALUE);
		LOOKUP_TABLE_K <= -- Make sure no index will fall out of boundary
			to_unsigned(0, 14) when IN_UNSIGNED <= 0 
		else
			to_unsigned(VECTOR_SIZE, 14) when IN_UNSIGNED >= VECTOR_SIZE 
		else
			IN_UNSIGNED;
  
		LOOKUP_TABLE_OUT <= TAN_SIG(to_integer(LOOKUP_TABLE_K));
		
		
		
		LOOKUP_TABLE_OUT_CONSTRAINED<=
			resize(LOOKUP_TABLE_OUT,U_SIZE,L_SIZE);
		

		UNIT_DELAY_PROCESS : process (clk)
			
			begin
				if CLK'event and CLK = '1' then
				UNIT_DELAY_OUT <= LOOKUP_TABLE_OUT_CONSTRAINED;
				end if;
		
		end process UNIT_DELAY_PROCESS;


		Y_VALUE <= UNIT_DELAY_OUT;
end RTL;
--=============================================================================
-- architecture end
--=============================================================================
